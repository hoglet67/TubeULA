module tube_ula(
      DACK
    , DRQ
    , HA0
    , HA1
    , HA2
    , HCS
    , HD0IN
    , HD0OUT
    , HD1IN
    , HD1OUT
    , HD2IN
    , HD2OUT
    , HD3IN
    , HD3OUT
    , HD4IN
    , HD4OUT
    , HD5IN
    , HD5OUT
    , HD6IN
    , HD6OUT
    , HD7IN
    , HD7OUT
    , HDOE
    , HIRQ
    , HO2
    , HRST
    , HRW
    , PA0
    , PA1
    , PA2
    , PCS
    , PD0IN
    , PD0OUT
    , PD1IN
    , PD1OUT
    , PD2IN
    , PD2OUT
    , PD3IN
    , PD3OUT
    , PD4IN
    , PD4OUT
    , PD5IN
    , PD5OUT
    , PD6IN
    , PD6OUT
    , PD7IN
    , PD7OUT
    , PDOE
    , PIRQ
    , PNMI
    , PNRDS
    , PNWDS
    , PRST
);
// Inputs
input DACK;
input HA0;
input HA1;
input HA2;
input HCS;
input HD0IN;
input HD1IN;
input HD2IN;
input HD3IN;
input HD4IN;
input HD5IN;
input HD6IN;
input HD7IN;
input HO2;
input HRST;
input HRW;
input PA0;
input PA1;
input PA2;
input PCS;
input PD0IN;
input PD1IN;
input PD2IN;
input PD3IN;
input PD4IN;
input PD5IN;
input PD6IN;
input PD7IN;
input PNRDS;
input PNWDS;
// Outputs
output DRQ;
output HD0OUT;
output HD1OUT;
output HD2OUT;
output HD3OUT;
output HD4OUT;
output HD5OUT;
output HD6OUT;
output HD7OUT;
output HDOE;
output HIRQ;
output PD0OUT;
output PD1OUT;
output PD2OUT;
output PD3OUT;
output PD4OUT;
output PD5OUT;
output PD6OUT;
output PD7OUT;
output PDOE;
output PIRQ;
output PNMI;
output PRST;
// Wires
wire HDOEA;
wire N1002;
wire N1003;
wire N1004;
wire N1035;
wire N1036;
wire N1037;
wire N1038;
wire N1039;
wire N1040;
wire N1041;
wire N1042;
wire N1043;
wire N1044;
wire N1046;
wire N1047;
wire N1048;
wire N1049;
wire N1050;
wire N1051;
wire N1052;
wire N1053;
wire N1056;
wire N1057;
wire N1058;
wire N1059;
wire N1060;
wire N1061;
wire N1062;
wire N1063;
wire N1064;
wire N1065;
wire N1066;
wire N1067;
wire N1068;
wire N1069;
wire N1070;
wire N1071;
wire N1072;
wire N1073;
wire N1074;
wire N1075;
wire N1076;
wire N1077;
wire N1078;
wire N1079;
wire N1080;
wire N1081;
wire N1082;
wire N1083;
wire N1084;
wire N1085;
wire N1086;
wire N1087;
wire N1089;
wire N1091;
wire N1093;
wire N1095;
wire N1097;
wire N1115;
wire N1117;
wire N1119;
wire N1121;
wire N1123;
wire N1125;
wire N1126;
wire N115;
wire N1155;
wire N116;
wire N117;
wire N118;
wire N1187;
wire N1188;
wire N1189;
wire N119;
wire N1190;
wire N1191;
wire N1192;
wire N1193;
wire N1194;
wire N1195;
wire N1196;
wire N1197;
wire N1198;
wire N1199;
wire N120;
wire N1200;
wire N1201;
wire N1202;
wire N1203;
wire N1204;
wire N1205;
wire N1206;
wire N1208;
wire N1209;
wire N121;
wire N1210;
wire N1211;
wire N1212;
wire N1213;
wire N1214;
wire N1215;
wire N1216;
wire N122;
wire N1226;
wire N1229;
wire N123;
wire N1232;
wire N1235;
wire N1238;
wire N124;
wire N1241;
wire N1244;
wire N1247;
wire N125;
wire N126;
wire N127;
wire N1313;
wire N1314;
wire N1315;
wire N1316;
wire N1317;
wire N1318;
wire N1319;
wire N1320;
wire N1321;
wire N1326;
wire N1327;
wire N1328;
wire N1329;
wire N1332;
wire N1335;
wire N1336;
wire N1339;
wire N1343;
wire N1346;
wire N1349;
wire N1396;
wire N1398;
wire N1399;
wire N140;
wire N141;
wire N1430;
wire N1431;
wire N1432;
wire N1433;
wire N1434;
wire N1435;
wire N1436;
wire N1437;
wire N1438;
wire N1439;
wire N1440;
wire N1441;
wire N1442;
wire N1443;
wire N1444;
wire N1445;
wire N1446;
wire N1447;
wire N1448;
wire N1449;
wire N1450;
wire N1451;
wire N1452;
wire N1453;
wire N1455;
wire N1456;
wire N1457;
wire N1458;
wire N1464;
wire N1466;
wire N1468;
wire N1470;
wire N1472;
wire N1474;
wire N1476;
wire N1478;
wire N1480;
wire N1482;
wire N1484;
wire N1486;
wire N1488;
wire N1490;
wire N1492;
wire N1494;
wire N1496;
wire N1498;
wire N1536;
wire N1537;
wire N1538;
wire N1570;
wire N1571;
wire N1572;
wire N1573;
wire N1574;
wire N1575;
wire N1576;
wire N1577;
wire N1578;
wire N1579;
wire N1580;
wire N1581;
wire N1582;
wire N1583;
wire N1584;
wire N1585;
wire N1586;
wire N1587;
wire N1588;
wire N1589;
wire N1590;
wire N1591;
wire N1592;
wire N1593;
wire N1594;
wire N1595;
wire N1596;
wire N1597;
wire N1598;
wire N1599;
wire N1600;
wire N1601;
wire N1602;
wire N1603;
wire N1604;
wire N1605;
wire N1606;
wire N1607;
wire N1608;
wire N1609;
wire N1610;
wire N1611;
wire N1612;
wire N1613;
wire N1614;
wire N1616;
wire N1617;
wire N1618;
wire N1619;
wire N1620;
wire N1622;
wire N1624;
wire N1626;
wire N1628;
wire N1630;
wire N1649;
wire N1651;
wire N1653;
wire N1655;
wire N1657;
wire N1687;
wire N1688;
wire N1719;
wire N1720;
wire N1721;
wire N1722;
wire N1723;
wire N1724;
wire N1725;
wire N1726;
wire N1727;
wire N1728;
wire N1729;
wire N1730;
wire N1731;
wire N1732;
wire N1733;
wire N1734;
wire N1735;
wire N1736;
wire N1737;
wire N1738;
wire N1739;
wire N1740;
wire N1741;
wire N1742;
wire N1743;
wire N1744;
wire N1745;
wire N1746;
wire N1748;
wire N175;
wire N1750;
wire N1759;
wire N176;
wire N1762;
wire N1765;
wire N1768;
wire N177;
wire N1771;
wire N1774;
wire N1777;
wire N1780;
wire N1817;
wire N1848;
wire N1849;
wire N1850;
wire N1851;
wire N1852;
wire N1853;
wire N1854;
wire N1855;
wire N1856;
wire N1857;
wire N1858;
wire N1859;
wire N1860;
wire N1861;
wire N1862;
wire N1863;
wire N1864;
wire N1865;
wire N1866;
wire N1867;
wire N1868;
wire N1869;
wire N1870;
wire N1871;
wire N1872;
wire N1873;
wire N1874;
wire N1875;
wire N1876;
wire N1877;
wire N1879;
wire N1882;
wire N1884;
wire N1886;
wire N1888;
wire N1890;
wire N1892;
wire N1894;
wire N1896;
wire N1898;
wire N1900;
wire N1902;
wire N1904;
wire N1906;
wire N1908;
wire N1910;
wire N1912;
wire N1914;
wire N1916;
wire N1955;
wire N1956;
wire N1988;
wire N1989;
wire N1990;
wire N1991;
wire N1992;
wire N1993;
wire N1994;
wire N1995;
wire N1996;
wire N1997;
wire N1998;
wire N1999;
wire N2000;
wire N2001;
wire N2002;
wire N2003;
wire N2004;
wire N2005;
wire N2006;
wire N2007;
wire N2008;
wire N2009;
wire N2010;
wire N2011;
wire N2012;
wire N2013;
wire N2014;
wire N2015;
wire N2016;
wire N2017;
wire N2018;
wire N2019;
wire N2020;
wire N2021;
wire N2022;
wire N2023;
wire N2024;
wire N2025;
wire N2026;
wire N2027;
wire N2028;
wire N2029;
wire N2030;
wire N2031;
wire N2032;
wire N2033;
wire N2034;
wire N2035;
wire N2036;
wire N2037;
wire N2038;
wire N2039;
wire N2040;
wire N2042;
wire N2044;
wire N2046;
wire N2048;
wire N2050;
wire N2069;
wire N207;
wire N2071;
wire N2073;
wire N2075;
wire N2077;
wire N2079;
wire N208;
wire N209;
wire N210;
wire N211;
wire N212;
wire N213;
wire N214;
wire N2140;
wire N2141;
wire N2142;
wire N2143;
wire N2144;
wire N2145;
wire N2146;
wire N2147;
wire N2148;
wire N2149;
wire N215;
wire N2150;
wire N2151;
wire N2152;
wire N2153;
wire N2154;
wire N2155;
wire N2156;
wire N2157;
wire N2158;
wire N2159;
wire N216;
wire N2160;
wire N2161;
wire N2162;
wire N2163;
wire N2164;
wire N2165;
wire N2166;
wire N2167;
wire N2168;
wire N217;
wire N2172;
wire N218;
wire N2181;
wire N2184;
wire N2187;
wire N219;
wire N2190;
wire N2193;
wire N2196;
wire N2199;
wire N220;
wire N2202;
wire N221;
wire N222;
wire N223;
wire N2239;
wire N2271;
wire N2272;
wire N2273;
wire N2274;
wire N2275;
wire N2276;
wire N2277;
wire N2278;
wire N2279;
wire N228;
wire N2280;
wire N2281;
wire N2282;
wire N2283;
wire N2284;
wire N2285;
wire N2286;
wire N2287;
wire N2288;
wire N2289;
wire N2290;
wire N2291;
wire N2292;
wire N2293;
wire N2294;
wire N2295;
wire N2296;
wire N2298;
wire N2299;
wire N23;
wire N230;
wire N2300;
wire N2301;
wire N2303;
wire N2306;
wire N2308;
wire N231;
wire N2310;
wire N2312;
wire N2314;
wire N2316;
wire N2318;
wire N2320;
wire N2322;
wire N2324;
wire N2326;
wire N2328;
wire N2330;
wire N2332;
wire N2334;
wire N2336;
wire N2338;
wire N234;
wire N2340;
wire N235;
wire N237;
wire N2379;
wire N2380;
wire N24;
wire N2412;
wire N2414;
wire N2415;
wire N2416;
wire N2417;
wire N2418;
wire N2419;
wire N2420;
wire N2421;
wire N2422;
wire N2423;
wire N2424;
wire N2425;
wire N2426;
wire N2427;
wire N2428;
wire N2429;
wire N2430;
wire N2431;
wire N2432;
wire N2433;
wire N2434;
wire N2435;
wire N2436;
wire N2437;
wire N2438;
wire N2439;
wire N2440;
wire N2441;
wire N2442;
wire N2443;
wire N2444;
wire N2445;
wire N2446;
wire N2447;
wire N2448;
wire N2449;
wire N2450;
wire N2451;
wire N2452;
wire N2453;
wire N2454;
wire N2455;
wire N2456;
wire N2457;
wire N2458;
wire N2459;
wire N2460;
wire N2461;
wire N2462;
wire N2463;
wire N2464;
wire N2465;
wire N2467;
wire N2469;
wire N2471;
wire N2473;
wire N2475;
wire N2494;
wire N2496;
wire N2498;
wire N25;
wire N2500;
wire N2502;
wire N2504;
wire N256;
wire N2565;
wire N2566;
wire N2567;
wire N2568;
wire N2569;
wire N2570;
wire N2571;
wire N2572;
wire N2573;
wire N2574;
wire N2575;
wire N2576;
wire N2577;
wire N2578;
wire N2579;
wire N2580;
wire N2581;
wire N2583;
wire N2584;
wire N2585;
wire N2586;
wire N2587;
wire N2588;
wire N2589;
wire N2590;
wire N2591;
wire N2592;
wire N2593;
wire N2594;
wire N2598;
wire N26;
wire N2607;
wire N2610;
wire N2613;
wire N2616;
wire N2619;
wire N2622;
wire N2625;
wire N2628;
wire N265;
wire N2665;
wire N269;
wire N2696;
wire N2697;
wire N2698;
wire N2699;
wire N27;
wire N2700;
wire N2701;
wire N2702;
wire N2703;
wire N2704;
wire N2705;
wire N2706;
wire N2707;
wire N2708;
wire N2709;
wire N2710;
wire N2711;
wire N2712;
wire N2713;
wire N2714;
wire N2715;
wire N2716;
wire N2717;
wire N2718;
wire N2719;
wire N2720;
wire N2721;
wire N2722;
wire N2723;
wire N2724;
wire N2725;
wire N2726;
wire N2729;
wire N2732;
wire N2734;
wire N2736;
wire N2738;
wire N2740;
wire N2742;
wire N2744;
wire N2746;
wire N2748;
wire N2750;
wire N2752;
wire N2754;
wire N2756;
wire N2758;
wire N2760;
wire N2762;
wire N2764;
wire N2766;
wire N28;
wire N2837;
wire N2838;
wire N2839;
wire N2840;
wire N2841;
wire N2842;
wire N2843;
wire N2844;
wire N2845;
wire N2846;
wire N2847;
wire N2848;
wire N2849;
wire N285;
wire N2850;
wire N2851;
wire N2852;
wire N2853;
wire N2854;
wire N2855;
wire N2856;
wire N2857;
wire N2859;
wire N286;
wire N2861;
wire N2862;
wire N2863;
wire N2864;
wire N2865;
wire N2866;
wire N2867;
wire N2868;
wire N2869;
wire N287;
wire N2870;
wire N2871;
wire N2872;
wire N2873;
wire N2874;
wire N2875;
wire N2876;
wire N2877;
wire N2878;
wire N2879;
wire N2880;
wire N2881;
wire N2882;
wire N2883;
wire N2884;
wire N2885;
wire N2887;
wire N2888;
wire N2889;
wire N2890;
wire N2891;
wire N2892;
wire N2894;
wire N2896;
wire N2898;
wire N2900;
wire N2902;
wire N2904;
wire N2923;
wire N2925;
wire N2927;
wire N2929;
wire N2931;
wire N2933;
wire N2993;
wire N2994;
wire N2995;
wire N2996;
wire N2997;
wire N2998;
wire N2999;
wire N3000;
wire N3001;
wire N3002;
wire N3003;
wire N3004;
wire N3005;
wire N3006;
wire N3007;
wire N3008;
wire N3009;
wire N3010;
wire N3011;
wire N3012;
wire N3013;
wire N3014;
wire N3015;
wire N3016;
wire N3017;
wire N3018;
wire N3019;
wire N3020;
wire N3021;
wire N3023;
wire N3033;
wire N3036;
wire N3039;
wire N3042;
wire N3045;
wire N3048;
wire N3051;
wire N3054;
wire N3093;
wire N31;
wire N3124;
wire N3125;
wire N3126;
wire N3127;
wire N3128;
wire N3129;
wire N3130;
wire N3131;
wire N3132;
wire N3133;
wire N3134;
wire N3135;
wire N3136;
wire N3137;
wire N3138;
wire N3139;
wire N3140;
wire N3141;
wire N3142;
wire N3143;
wire N3144;
wire N3145;
wire N3146;
wire N3147;
wire N3148;
wire N3149;
wire N3150;
wire N3151;
wire N3153;
wire N3154;
wire N3156;
wire N3157;
wire N3158;
wire N3160;
wire N3164;
wire N3166;
wire N3168;
wire N317;
wire N3170;
wire N3172;
wire N3174;
wire N3176;
wire N3178;
wire N318;
wire N3180;
wire N3182;
wire N3184;
wire N3186;
wire N3188;
wire N319;
wire N3190;
wire N3192;
wire N3194;
wire N3196;
wire N3198;
wire N32;
wire N320;
wire N3200;
wire N321;
wire N322;
wire N323;
wire N3237;
wire N3238;
wire N324;
wire N325;
wire N326;
wire N327;
wire N3270;
wire N3271;
wire N3272;
wire N3273;
wire N3274;
wire N3275;
wire N3276;
wire N3277;
wire N3278;
wire N3279;
wire N328;
wire N3280;
wire N3281;
wire N3282;
wire N3283;
wire N3284;
wire N3285;
wire N3286;
wire N3287;
wire N3288;
wire N3289;
wire N329;
wire N3291;
wire N3292;
wire N3293;
wire N3294;
wire N3295;
wire N3296;
wire N3297;
wire N3298;
wire N3299;
wire N33;
wire N330;
wire N3300;
wire N3301;
wire N3302;
wire N3303;
wire N3304;
wire N3305;
wire N3306;
wire N3307;
wire N3308;
wire N3309;
wire N331;
wire N3310;
wire N3311;
wire N3312;
wire N3313;
wire N3314;
wire N3315;
wire N3316;
wire N3317;
wire N3318;
wire N3319;
wire N332;
wire N3320;
wire N3321;
wire N3322;
wire N3323;
wire N3325;
wire N3327;
wire N3329;
wire N333;
wire N3331;
wire N3333;
wire N334;
wire N335;
wire N3352;
wire N3354;
wire N3356;
wire N3358;
wire N3360;
wire N3362;
wire N338;
wire N34;
wire N3423;
wire N3424;
wire N3425;
wire N3426;
wire N3427;
wire N3428;
wire N3429;
wire N343;
wire N3430;
wire N3431;
wire N3432;
wire N3433;
wire N3434;
wire N3435;
wire N3436;
wire N3437;
wire N3438;
wire N3439;
wire N3440;
wire N3441;
wire N3442;
wire N3443;
wire N3444;
wire N3445;
wire N3446;
wire N3447;
wire N3448;
wire N3449;
wire N3450;
wire N3451;
wire N3455;
wire N3464;
wire N3467;
wire N347;
wire N3470;
wire N3473;
wire N3476;
wire N3479;
wire N3482;
wire N3485;
wire N35;
wire N350;
wire N3522;
wire N3554;
wire N3555;
wire N3556;
wire N3557;
wire N3558;
wire N3559;
wire N3560;
wire N3561;
wire N3562;
wire N3563;
wire N3564;
wire N3565;
wire N3566;
wire N3567;
wire N3568;
wire N3569;
wire N3570;
wire N3571;
wire N3572;
wire N3573;
wire N3574;
wire N3575;
wire N3576;
wire N3577;
wire N3578;
wire N3579;
wire N3580;
wire N3582;
wire N3583;
wire N3584;
wire N3585;
wire N3587;
wire N3590;
wire N3592;
wire N3594;
wire N3596;
wire N3598;
wire N36;
wire N3600;
wire N3602;
wire N3604;
wire N3606;
wire N3608;
wire N3610;
wire N3612;
wire N3614;
wire N3616;
wire N3618;
wire N3620;
wire N3622;
wire N3624;
wire N3626;
wire N364;
wire N3664;
wire N3665;
wire N3697;
wire N3698;
wire N3699;
wire N37;
wire N3700;
wire N3701;
wire N3702;
wire N3703;
wire N3704;
wire N3705;
wire N3706;
wire N3707;
wire N3708;
wire N3709;
wire N3710;
wire N3711;
wire N3712;
wire N3713;
wire N3714;
wire N3715;
wire N3716;
wire N3718;
wire N3719;
wire N372;
wire N3720;
wire N3721;
wire N3722;
wire N3723;
wire N3724;
wire N3725;
wire N3726;
wire N3727;
wire N3728;
wire N3729;
wire N3730;
wire N3731;
wire N3732;
wire N3733;
wire N3734;
wire N3735;
wire N3736;
wire N3737;
wire N3738;
wire N3739;
wire N3740;
wire N3741;
wire N3742;
wire N3743;
wire N3744;
wire N3745;
wire N3746;
wire N3747;
wire N3748;
wire N3749;
wire N3750;
wire N3752;
wire N3754;
wire N3756;
wire N3758;
wire N3760;
wire N3779;
wire N3781;
wire N3783;
wire N3785;
wire N3787;
wire N3789;
wire N38;
wire N384;
wire N3851;
wire N3852;
wire N3853;
wire N3854;
wire N3855;
wire N3856;
wire N3857;
wire N3858;
wire N3859;
wire N3860;
wire N3861;
wire N3862;
wire N3863;
wire N3864;
wire N3865;
wire N3866;
wire N3867;
wire N3868;
wire N3869;
wire N3870;
wire N3871;
wire N3872;
wire N3873;
wire N3874;
wire N3875;
wire N3876;
wire N3877;
wire N3878;
wire N3879;
wire N3883;
wire N3892;
wire N3895;
wire N3898;
wire N39;
wire N390;
wire N3901;
wire N3904;
wire N3907;
wire N3910;
wire N3913;
wire N3950;
wire N397;
wire N398;
wire N3982;
wire N3983;
wire N3984;
wire N3985;
wire N3986;
wire N3987;
wire N3988;
wire N3989;
wire N399;
wire N3990;
wire N3991;
wire N3992;
wire N3993;
wire N3994;
wire N3995;
wire N3996;
wire N3997;
wire N3998;
wire N3999;
wire N40;
wire N4000;
wire N4001;
wire N4002;
wire N4003;
wire N4004;
wire N4005;
wire N4006;
wire N4007;
wire N4009;
wire N4010;
wire N4011;
wire N4012;
wire N4014;
wire N4017;
wire N4019;
wire N4021;
wire N4023;
wire N4025;
wire N4027;
wire N4029;
wire N4031;
wire N4033;
wire N4035;
wire N4037;
wire N4039;
wire N4041;
wire N4043;
wire N4045;
wire N4047;
wire N4049;
wire N4051;
wire N4090;
wire N4091;
wire N4123;
wire N4124;
wire N4125;
wire N4126;
wire N4127;
wire N4128;
wire N4129;
wire N4130;
wire N4131;
wire N4132;
wire N4133;
wire N4134;
wire N4135;
wire N4136;
wire N4137;
wire N4138;
wire N4139;
wire N4140;
wire N4141;
wire N4142;
wire N4144;
wire N4145;
wire N4146;
wire N4147;
wire N4148;
wire N4149;
wire N4150;
wire N4151;
wire N4152;
wire N4153;
wire N4154;
wire N4155;
wire N4156;
wire N4157;
wire N4158;
wire N4159;
wire N4160;
wire N4161;
wire N4162;
wire N4163;
wire N4164;
wire N4165;
wire N4166;
wire N4167;
wire N4168;
wire N4169;
wire N4170;
wire N4171;
wire N4172;
wire N4173;
wire N4174;
wire N4175;
wire N4176;
wire N4178;
wire N4180;
wire N4182;
wire N4184;
wire N4186;
wire N4205;
wire N4207;
wire N4209;
wire N4211;
wire N4213;
wire N4215;
wire N4276;
wire N4277;
wire N4278;
wire N4279;
wire N4280;
wire N4281;
wire N4282;
wire N4283;
wire N4284;
wire N4285;
wire N4286;
wire N4287;
wire N4288;
wire N4289;
wire N4290;
wire N4291;
wire N4292;
wire N4293;
wire N4294;
wire N4295;
wire N4296;
wire N4297;
wire N4298;
wire N4299;
wire N430;
wire N4300;
wire N4301;
wire N4302;
wire N4303;
wire N4304;
wire N4307;
wire N431;
wire N4316;
wire N4319;
wire N432;
wire N4322;
wire N4325;
wire N4328;
wire N433;
wire N4331;
wire N4334;
wire N4337;
wire N434;
wire N435;
wire N436;
wire N437;
wire N4375;
wire N438;
wire N439;
wire N440;
wire N4406;
wire N4407;
wire N4408;
wire N4409;
wire N441;
wire N4410;
wire N4411;
wire N4412;
wire N4413;
wire N442;
wire N443;
wire N444;
wire N445;
wire N446;
wire N447;
wire N448;
wire N449;
wire N450;
wire N451;
wire N452;
wire N453;
wire N454;
wire N455;
wire N456;
wire N457;
wire N459;
wire N462;
wire N464;
wire N466;
wire N468;
wire N470;
wire N472;
wire N473;
wire N475;
wire N476;
wire N478;
wire N479;
wire N481;
wire N483;
wire N486;
wire N488;
wire N490;
wire N492;
wire N493;
wire N496;
wire N498;
wire N50;
wire N507;
wire N510;
wire N514;
wire N518;
wire N522;
wire N526;
wire N530;
wire N533;
wire N541;
wire N542;
wire N543;
wire N544;
wire N545;
wire N546;
wire N547;
wire N578;
wire N579;
wire N580;
wire N581;
wire N582;
wire N583;
wire N584;
wire N585;
wire N586;
wire N587;
wire N588;
wire N589;
wire N590;
wire N591;
wire N592;
wire N594;
wire N595;
wire N596;
wire N597;
wire N598;
wire N599;
wire N600;
wire N601;
wire N602;
wire N603;
wire N604;
wire N628;
wire N632;
wire N638;
wire N641;
wire N644;
wire N647;
wire N650;
wire N653;
wire N656;
wire N659;
wire N662;
wire N664;
wire N666;
wire N701;
wire N702;
wire N703;
wire N704;
wire N705;
wire N706;
wire N707;
wire N708;
wire N709;
wire N710;
wire N711;
wire N712;
wire N713;
wire N714;
wire N715;
wire N716;
wire N717;
wire N718;
wire N719;
wire N720;
wire N721;
wire N722;
wire N723;
wire N724;
wire N725;
wire N737;
wire N772;
wire N792;
wire N799;
wire N800;
wire N801;
wire N802;
wire N803;
wire N804;
wire N805;
wire N806;
wire N807;
wire N808;
wire N809;
wire N818;
wire N819;
wire N822;
wire N823;
wire N824;
wire N825;
wire N826;
wire N827;
wire N828;
wire N829;
wire N830;
wire N831;
wire N832;
wire N833;
wire N834;
wire N835;
wire N837;
wire N839;
wire N84;
wire N876;
wire N899;
wire N900;
wire N901;
wire N902;
wire N903;
wire N904;
wire N905;
wire N906;
wire N907;
wire N908;
wire N909;
wire N910;
wire N911;
wire N912;
wire N913;
wire N914;
wire N915;
wire N916;
wire N917;
wire N918;
wire N919;
wire N920;
wire N921;
wire N922;
wire N923;
wire N924;
wire N926;
wire N932;
wire N934;
wire N936;
wire N938;
wire N940;
wire N942;
wire N944;
wire N946;
wire N948;
wire N950;
wire N952;
wire N954;
wire N956;
wire N958;
wire N960;
wire N962;
wire N967;
wire N974;
wire PDOEA;
wire PDOEB;
wire _HD0IN;
wire _HD1IN;
wire _HD2IN;
wire _HD3IN;
wire _HD4IN;
wire _HD5IN;
wire _HD6IN;
wire _HD7IN;
nor #5 GDRQ(DRQ,N321);
nor #5 GHD0OUT(HD0OUT,N4007,N4012,N4142,N4175,N4215);
nor #5 GHD1OUT(HD1OUT,N3580,N3585,N3716,N3749,N3789);
nor #5 GHD2OUT(HD2OUT,N3151,N3158,N3289,N3322,N3362);
nor #5 GHD3OUT(HD3OUT,N2725,N2726,N2856,N2857,N2933);
nor #5 GHD4OUT(HD4OUT,N2296,N2301,N2432,N2464,N2504);
nor #5 GHD5OUT(HD5OUT,N1873,N1877,N2007,N2039,N2079);
nor #5 GHD6OUT(HD6OUT,N1335,N1336,N1436,N1437,N1458,N1588,N1620,N1687);
nor #5 GHD7OUT(HD7OUT,N1035,N1083,N1125,N1155,N1187,N899,N921,N967);
nor #5 GHDOEA(HDOEA,HCS,N116,N50);
nor #5 GHIRQ(HIRQ,N1432);
nor #5 GN1002(N1002,N1060,N1093);
nor #5 GN1003(N1003,N903);
nor #5 GN1004(N1004,N1080,N1117);
nor #5 GN1035(N1035,N1004,N441);
nor #5 GN1036(N1036,N1057,N459);
nor #5 GN1037(N1037,N701,N934);
nor #5 GN1038(N1038,N702,N938);
nor #5 GN1039(N1039,N703,N942);
nor #5 GN1040(N1040,N704,N946);
nor #5 GN1041(N1041,N705,N950);
nor #5 GN1042(N1042,N706,N954);
nor #5 GN1043(N1043,N707,N958);
nor #5 GN1044(N1044,N1201,N792);
nor #5 GN1046(N1046,N601,N904);
nor #5 GN1047(N1047,N510,N906);
nor #5 GN1048(N1048,N579,N908);
nor #5 GN1049(N1049,N581,N910);
nor #5 GN1050(N1050,N583,N912);
nor #5 GN1051(N1051,N585,N914);
nor #5 GN1052(N1052,N587,N916);
nor #5 GN1053(N1053,N589,N918);
nor #5 GN1056(N1056,N34,N709);
nor #5 GN1057(N1057,N1059,N1091);
nor #5 GN1058(N1058,N1084,N1189);
nor #5 GN1059(N1059,N1057,N1190);
nor #5 GN1060(N1060,N1002,N1191);
nor #5 GN1061(N1061,N1192,N923);
nor #5 GN1062(N1062,N1085,N1193);
nor #5 GN1063(N1063,N1064,N904);
nor #5 GN1064(N1064,N1046,N1063);
nor #5 GN1065(N1065,N1066,N906);
nor #5 GN1066(N1066,N1047,N1065);
nor #5 GN1067(N1067,N1068,N908);
nor #5 GN1068(N1068,N1048,N1067);
nor #5 GN1069(N1069,N1070,N910);
nor #5 GN1070(N1070,N1049,N1069);
nor #5 GN1071(N1071,N1072,N912);
nor #5 GN1072(N1072,N1050,N1071);
nor #5 GN1073(N1073,N1074,N914);
nor #5 GN1074(N1074,N1051,N1073);
nor #5 GN1075(N1075,N1076,N916);
nor #5 GN1076(N1076,N1052,N1075);
nor #5 GN1077(N1077,N1078,N918);
nor #5 GN1078(N1078,N1053,N1077);
nor #5 GN1079(N1079,N1086,N1202);
nor #5 GN1080(N1080,N1004,N1203);
nor #5 GN1081(N1081,N1204,N920);
nor #5 GN1082(N1082,N1121,N1123);
nor #5 GN1083(N1083,N37,N664);
nor #5 GN1084(N1084,N1058,N1089);
nor #5 GN1085(N1085,N1062,N1097);
nor #5 GN1086(N1086,N1079,N1115);
nor #5 GN1087(N1087,N120,N628);
nor #5 GN1089(N1089,N710,N824);
nor #5 GN1091(N1091,N1190,N808);
nor #5 GN1093(N1093,N1191,N809);
nor #5 GN1095(N1095,N1192,N632);
nor #5 GN1097(N1097,N1193,N338);
nor #5 GN1115(N1115,N1202,N835);
nor #5 GN1117(N1117,N1203,N662);
nor #5 GN1119(N1119,N1204,N818);
nor #5 GN1121(N1121,N1082,N1205);
nor #5 GN1123(N1123,N1205,N819);
nor #5 GN1125(N1125,N498,N919);
nor #5 GN1126(N1126,N1058,N442);
nor #5 GN115(N115,N124,N35);
nor #5 GN1155(N1155,N343,N84);
nor #5 GN116(N116,HO2);
nor #5 GN117(N117,N122);
nor #5 GN118(N118,N24);
nor #5 GN1187(N1187,N1082,N334);
nor #5 GN1188(N1188,N118,N1208);
nor #5 GN1189(N1189,N1089,N824);
nor #5 GN119(N119,N36);
nor #5 GN1190(N1190,N710,N808);
nor #5 GN1191(N1191,N710,N809);
nor #5 GN1192(N1192,N1062,N632);
nor #5 GN1193(N1193,N338,N710);
nor #5 GN1194(N1194,N1209,N1226);
nor #5 GN1195(N1195,N1210,N1229);
nor #5 GN1196(N1196,N1211,N1232);
nor #5 GN1197(N1197,N1212,N1235);
nor #5 GN1198(N1198,N1213,N1238);
nor #5 GN1199(N1199,N1214,N1241);
nor #5 GN120(N120,N123);
nor #5 GN1200(N1200,N1215,N1244);
nor #5 GN1201(N1201,N1216,N1247);
nor #5 GN1202(N1202,N823,N835);
nor #5 GN1203(N1203,N1079,N662);
nor #5 GN1204(N1204,N818,N823);
nor #5 GN1205(N1205,N819,N823);
nor #5 GN1206(N1206,N332,N595);
nor #5 GN1208(N1208,N321);
nor #5 GN1209(N1209,N1063,N800);
nor #5 GN121(N121,HCS,N116,N50);
nor #5 GN1210(N1210,N1065,N801);
nor #5 GN1211(N1211,N1067,N802);
nor #5 GN1212(N1212,N1069,N803);
nor #5 GN1213(N1213,N1071,N804);
nor #5 GN1214(N1214,N1073,N805);
nor #5 GN1215(N1215,N1075,N806);
nor #5 GN1216(N1216,N1077,N807);
nor #5 GN122(N122,HA0,HA2,N39);
nor #5 GN1226(N1226,N1194,N1313);
nor #5 GN1229(N1229,N1195,N1315);
nor #5 GN123(N123,N23,N32,PA0,PA2);
nor #5 GN1232(N1232,N1196,N1316);
nor #5 GN1235(N1235,N1197,N1317);
nor #5 GN1238(N1238,N1198,N1318);
nor #5 GN124(N124,PCS,PNWDS);
nor #5 GN1241(N1241,N1199,N1319);
nor #5 GN1244(N1244,N1200,N1320);
nor #5 GN1247(N1247,N1201,N1321);
nor #5 GN125(N125,N126,N176);
nor #5 GN126(N126,PCS,PNRDS);
nor #5 GN127(N127,N121);
nor #5 GN1313(N1313,N1209,N800);
nor #5 GN1314(N1314,N664);
nor #5 GN1315(N1315,N1210,N801);
nor #5 GN1316(N1316,N1211,N802);
nor #5 GN1317(N1317,N1212,N803);
nor #5 GN1318(N1318,N1213,N804);
nor #5 GN1319(N1319,N1214,N805);
nor #5 GN1320(N1320,N1215,N806);
nor #5 GN1321(N1321,N1216,N807);
nor #5 GN1326(N1326,N1346);
nor #5 GN1327(N1327,N708);
nor #5 GN1328(N1328,N1314,N34);
nor #5 GN1329(N1329,N118,N1339);
nor #5 GN1332(N1332,N1343,N321);
nor #5 GN1335(N1335,N318,N84);
nor #5 GN1336(N1336,N1327,N335);
nor #5 GN1339(N1339,N343);
nor #5 GN1343(N1343,N1434);
nor #5 GN1346(N1346,N4011,N4017,N4123);
nor #5 GN1349(N1349,N1617,N1719);
nor #5 GN1396(N1396,N1496,N1498);
nor #5 GN1398(N1398,N120,N1430);
nor #5 GN1399(N1399,N628);
nor #5 GN140(N140,N23,PA0,PA1,PA2);
nor #5 GN141(N141,HA0,HA1,HA2);
nor #5 GN1430(N1430,N666);
nor #5 GN1431(N1431,N1736,N1750);
nor #5 GN1432(N1432,N1314,N1326);
nor #5 GN1433(N1433,N1876,N1882,N1988);
nor #5 GN1434(N1434,N2724,N2732,N2837);
nor #5 GN1435(N1435,N1349,N442);
nor #5 GN1436(N1436,N117,N1399);
nor #5 GN1437(N1437,N1396,N498);
nor #5 GN1438(N1438,N1431,N601);
nor #5 GN1439(N1439,N1468,N1470);
nor #5 GN1440(N1440,N1439,N510);
nor #5 GN1441(N1441,N1472,N1474);
nor #5 GN1442(N1442,N1441,N579);
nor #5 GN1443(N1443,N1476,N1478);
nor #5 GN1444(N1444,N1443,N581);
nor #5 GN1445(N1445,N1480,N1482);
nor #5 GN1446(N1446,N1445,N583);
nor #5 GN1447(N1447,N1484,N1486);
nor #5 GN1448(N1448,N1447,N585);
nor #5 GN1449(N1449,N1488,N1490);
nor #5 GN1450(N1450,N1449,N587);
nor #5 GN1451(N1451,N1492,N1494);
nor #5 GN1452(N1452,N1451,N589);
nor #5 GN1453(N1453,N709);
nor #5 GN1455(N1455,N325,N454);
nor #5 GN1456(N1456,N1592,N1628);
nor #5 GN1457(N1457,N1466,N435);
nor #5 GN1458(N1458,N1453,N37);
nor #5 GN1464(N1464,N1571,N924);
nor #5 GN1466(N1466,N1206,N1570,N1571);
nor #5 GN1468(N1468,N1439,N1572);
nor #5 GN1470(N1470,N1724,N701);
nor #5 GN1472(N1472,N1441,N1573);
nor #5 GN1474(N1474,N1725,N702);
nor #5 GN1476(N1476,N1443,N1574);
nor #5 GN1478(N1478,N1726,N703);
nor #5 GN1480(N1480,N1445,N1575);
nor #5 GN1482(N1482,N1727,N704);
nor #5 GN1484(N1484,N1447,N1576);
nor #5 GN1486(N1486,N1728,N705);
nor #5 GN1488(N1488,N1449,N1577);
nor #5 GN1490(N1490,N1729,N706);
nor #5 GN1492(N1492,N1451,N1578);
nor #5 GN1494(N1494,N1730,N707);
nor #5 GN1496(N1496,N1396,N1579);
nor #5 GN1498(N1498,N1579,N792);
nor #5 GN1536(N1536,N1456,N326);
nor #5 GN1537(N1537,N1591,N1626);
nor #5 GN1538(N1538,N1611,N1651);
nor #5 GN1570(N1570,N1206,N924);
nor #5 GN1571(N1571,N1745,N1746);
nor #5 GN1572(N1572,N1470,N701);
nor #5 GN1573(N1573,N1474,N702);
nor #5 GN1574(N1574,N1478,N703);
nor #5 GN1575(N1575,N1482,N704);
nor #5 GN1576(N1576,N1486,N705);
nor #5 GN1577(N1577,N1490,N706);
nor #5 GN1578(N1578,N1494,N707);
nor #5 GN1579(N1579,N1731,N792);
nor #5 GN1580(N1580,N1438,N601);
nor #5 GN1581(N1581,N1440,N510);
nor #5 GN1582(N1582,N1442,N579);
nor #5 GN1583(N1583,N1444,N581);
nor #5 GN1584(N1584,N1446,N583);
nor #5 GN1585(N1585,N1448,N585);
nor #5 GN1586(N1586,N1450,N587);
nor #5 GN1587(N1587,N1452,N589);
nor #5 GN1588(N1588,N1538,N441);
nor #5 GN1589(N1589,N1590,N1624);
nor #5 GN1590(N1590,N1589,N1720);
nor #5 GN1591(N1591,N1537,N1721);
nor #5 GN1592(N1592,N1456,N1722);
nor #5 GN1593(N1593,N1618,N1723);
nor #5 GN1594(N1594,N1438,N1595);
nor #5 GN1595(N1595,N1580,N1594);
nor #5 GN1596(N1596,N1440,N1597);
nor #5 GN1597(N1597,N1581,N1596);
nor #5 GN1598(N1598,N1442,N1599);
nor #5 GN1599(N1599,N1582,N1598);
nor #5 GN1600(N1600,N1444,N1601);
nor #5 GN1601(N1601,N1583,N1600);
nor #5 GN1602(N1602,N1446,N1603);
nor #5 GN1603(N1603,N1584,N1602);
nor #5 GN1604(N1604,N1448,N1605);
nor #5 GN1605(N1605,N1585,N1604);
nor #5 GN1606(N1606,N1450,N1607);
nor #5 GN1607(N1607,N1586,N1606);
nor #5 GN1608(N1608,N1452,N1609);
nor #5 GN1609(N1609,N1587,N1608);
nor #5 GN1610(N1610,N1619,N1732);
nor #5 GN1611(N1611,N1538,N1733);
nor #5 GN1612(N1612,N1613,N1653);
nor #5 GN1613(N1613,N1612,N1734);
nor #5 GN1614(N1614,N1655,N1657);
nor #5 GN1616(N1616,N1537,N327);
nor #5 GN1617(N1617,N1349,N1622);
nor #5 GN1618(N1618,N1593,N1630);
nor #5 GN1619(N1619,N1610,N1649);
nor #5 GN1620(N1620,N1612,N496);
nor #5 GN1622(N1622,N1571,N824);
nor #5 GN1624(N1624,N1720,N808);
nor #5 GN1626(N1626,N1721,N809);
nor #5 GN1628(N1628,N1722,N632);
nor #5 GN1630(N1630,N1723,N338);
nor #5 GN1649(N1649,N1732,N835);
nor #5 GN1651(N1651,N1733,N662);
nor #5 GN1653(N1653,N1734,N818);
nor #5 GN1655(N1655,N1614,N1735);
nor #5 GN1657(N1657,N1735,N819);
nor #5 GN1687(N1687,N1614,N334);
nor #5 GN1688(N1688,N1589,N459);
nor #5 GN1719(N1719,N1622,N824);
nor #5 GN1720(N1720,N1571,N808);
nor #5 GN1721(N1721,N1571,N809);
nor #5 GN1722(N1722,N1593,N632);
nor #5 GN1723(N1723,N1571,N338);
nor #5 GN1724(N1724,N1737,N1759);
nor #5 GN1725(N1725,N1738,N1762);
nor #5 GN1726(N1726,N1739,N1765);
nor #5 GN1727(N1727,N1740,N1768);
nor #5 GN1728(N1728,N1741,N1771);
nor #5 GN1729(N1729,N1742,N1774);
nor #5 GN1730(N1730,N1743,N1777);
nor #5 GN1731(N1731,N1744,N1780);
nor #5 GN1732(N1732,N1431,N835);
nor #5 GN1733(N1733,N1610,N662);
nor #5 GN1734(N1734,N1431,N818);
nor #5 GN1735(N1735,N1431,N819);
nor #5 GN1736(N1736,N115,N1748);
nor #5 GN1737(N1737,N1594,N800);
nor #5 GN1738(N1738,N1596,N801);
nor #5 GN1739(N1739,N1598,N802);
nor #5 GN1740(N1740,N1600,N803);
nor #5 GN1741(N1741,N1602,N804);
nor #5 GN1742(N1742,N1604,N805);
nor #5 GN1743(N1743,N1606,N806);
nor #5 GN1744(N1744,N1608,N807);
nor #5 GN1745(N1745,N1571,N1817);
nor #5 GN1746(N1746,N26,_HD6IN);
nor #5 GN1748(N1748,N115,PD6IN);
nor #5 GN175(N175,N124,N35);
nor #5 GN1750(N1750,N1431,N1748);
nor #5 GN1759(N1759,N1724,N1849);
nor #5 GN176(N176,DACK,PNWDS);
nor #5 GN1762(N1762,N1725,N1850);
nor #5 GN1765(N1765,N1726,N1851);
nor #5 GN1768(N1768,N1727,N1852);
nor #5 GN177(N177,N175,N459);
nor #5 GN1771(N1771,N1728,N1853);
nor #5 GN1774(N1774,N1729,N1854);
nor #5 GN1777(N1777,N1730,N1855);
nor #5 GN1780(N1780,N1731,N1856);
nor #5 GN1817(N1817,N1746,N26);
nor #5 GN1848(N1848,N2158,N2172);
nor #5 GN1849(N1849,N1737,N800);
nor #5 GN1850(N1850,N1738,N801);
nor #5 GN1851(N1851,N1739,N802);
nor #5 GN1852(N1852,N1740,N803);
nor #5 GN1853(N1853,N1741,N804);
nor #5 GN1854(N1854,N1742,N805);
nor #5 GN1855(N1855,N1743,N806);
nor #5 GN1856(N1856,N1744,N807);
nor #5 GN1857(N1857,N1848,N601);
nor #5 GN1858(N1858,N1886,N1888);
nor #5 GN1859(N1859,N1858,N510);
nor #5 GN1860(N1860,N1890,N1892);
nor #5 GN1861(N1861,N1860,N579);
nor #5 GN1862(N1862,N1894,N1896);
nor #5 GN1863(N1863,N1862,N581);
nor #5 GN1864(N1864,N1898,N1900);
nor #5 GN1865(N1865,N1864,N583);
nor #5 GN1866(N1866,N1902,N1904);
nor #5 GN1867(N1867,N1866,N585);
nor #5 GN1868(N1868,N1906,N1908);
nor #5 GN1869(N1869,N1868,N587);
nor #5 GN1870(N1870,N1910,N1912);
nor #5 GN1871(N1871,N1870,N589);
nor #5 GN1872(N1872,N1914,N1916);
nor #5 GN1873(N1873,N1433,N335);
nor #5 GN1874(N1874,N1433,N325);
nor #5 GN1875(N1875,N2013,N2048);
nor #5 GN1876(N1876,N1433,N1884);
nor #5 GN1877(N1877,N1872,N498);
nor #5 GN1879(N1879,N1875,N326);
nor #5 GN1882(N1882,N1990,N924);
nor #5 GN1884(N1884,N1206,N1988,N1990);
nor #5 GN1886(N1886,N1858,N1991);
nor #5 GN1888(N1888,N2145,N701);
nor #5 GN1890(N1890,N1860,N1992);
nor #5 GN1892(N1892,N2146,N702);
nor #5 GN1894(N1894,N1862,N1993);
nor #5 GN1896(N1896,N2147,N703);
nor #5 GN1898(N1898,N1864,N1994);
nor #5 GN1900(N1900,N2148,N704);
nor #5 GN1902(N1902,N1866,N1995);
nor #5 GN1904(N1904,N2149,N705);
nor #5 GN1906(N1906,N1868,N1996);
nor #5 GN1908(N1908,N2150,N706);
nor #5 GN1910(N1910,N1870,N1997);
nor #5 GN1912(N1912,N2151,N707);
nor #5 GN1914(N1914,N1872,N1998);
nor #5 GN1916(N1916,N1998,N792);
nor #5 GN1955(N1955,N2012,N2046);
nor #5 GN1956(N1956,N2032,N2071);
nor #5 GN1988(N1988,N1206,N924);
nor #5 GN1989(N1989,N1955,N327);
nor #5 GN1990(N1990,N2167,N2168);
nor #5 GN1991(N1991,N1888,N701);
nor #5 GN1992(N1992,N1892,N702);
nor #5 GN1993(N1993,N1896,N703);
nor #5 GN1994(N1994,N1900,N704);
nor #5 GN1995(N1995,N1904,N705);
nor #5 GN1996(N1996,N1908,N706);
nor #5 GN1997(N1997,N1912,N707);
nor #5 GN1998(N1998,N2152,N792);
nor #5 GN1999(N1999,N1857,N601);
nor #5 GN2000(N2000,N1859,N510);
nor #5 GN2001(N2001,N1861,N579);
nor #5 GN2002(N2002,N1863,N581);
nor #5 GN2003(N2003,N1865,N583);
nor #5 GN2004(N2004,N1867,N585);
nor #5 GN2005(N2005,N1869,N587);
nor #5 GN2006(N2006,N1871,N589);
nor #5 GN2007(N2007,N1956,N441);
nor #5 GN2008(N2008,N2010,N442);
nor #5 GN2009(N2009,N2011,N2044);
nor #5 GN2010(N2010,N2036,N2140);
nor #5 GN2011(N2011,N2009,N2141);
nor #5 GN2012(N2012,N1955,N2142);
nor #5 GN2013(N2013,N1875,N2143);
nor #5 GN2014(N2014,N2037,N2144);
nor #5 GN2015(N2015,N1857,N2016);
nor #5 GN2016(N2016,N1999,N2015);
nor #5 GN2017(N2017,N1859,N2018);
nor #5 GN2018(N2018,N2000,N2017);
nor #5 GN2019(N2019,N1861,N2020);
nor #5 GN2020(N2020,N2001,N2019);
nor #5 GN2021(N2021,N1863,N2022);
nor #5 GN2022(N2022,N2002,N2021);
nor #5 GN2023(N2023,N1865,N2024);
nor #5 GN2024(N2024,N2003,N2023);
nor #5 GN2025(N2025,N1867,N2026);
nor #5 GN2026(N2026,N2004,N2025);
nor #5 GN2027(N2027,N1869,N2028);
nor #5 GN2028(N2028,N2005,N2027);
nor #5 GN2029(N2029,N1871,N2030);
nor #5 GN2030(N2030,N2006,N2029);
nor #5 GN2031(N2031,N2038,N2153);
nor #5 GN2032(N2032,N1956,N2154);
nor #5 GN2033(N2033,N2034,N2073);
nor #5 GN2034(N2034,N2033,N2155);
nor #5 GN2035(N2035,N2075,N2077);
nor #5 GN2036(N2036,N2010,N2042);
nor #5 GN2037(N2037,N2014,N2050);
nor #5 GN2038(N2038,N2031,N2069);
nor #5 GN2039(N2039,N2033,N496);
nor #5 GN2040(N2040,N2009,N459);
nor #5 GN2042(N2042,N1990,N824);
nor #5 GN2044(N2044,N2141,N808);
nor #5 GN2046(N2046,N2142,N809);
nor #5 GN2048(N2048,N2143,N632);
nor #5 GN2050(N2050,N2144,N338);
nor #5 GN2069(N2069,N2153,N835);
nor #5 GN207(N207,N119,N498);
nor #5 GN2071(N2071,N2154,N662);
nor #5 GN2073(N2073,N2155,N818);
nor #5 GN2075(N2075,N2035,N2156);
nor #5 GN2077(N2077,N2156,N819);
nor #5 GN2079(N2079,N2035,N334);
nor #5 GN208(N208,N119,N496);
nor #5 GN209(N209,N175,N327);
nor #5 GN210(N210,N235,N237);
nor #5 GN211(N211,N23,N31,PA1,PA2);
nor #5 GN212(N212,N23,N31,N32,PA2);
nor #5 GN213(N213,N31,N33,PA1);
nor #5 GN214(N214,N23,N31,N32,N33);
nor #5 GN2140(N2140,N2042,N824);
nor #5 GN2141(N2141,N1990,N808);
nor #5 GN2142(N2142,N1990,N809);
nor #5 GN2143(N2143,N2014,N632);
nor #5 GN2144(N2144,N1990,N338);
nor #5 GN2145(N2145,N2159,N2181);
nor #5 GN2146(N2146,N2160,N2184);
nor #5 GN2147(N2147,N2161,N2187);
nor #5 GN2148(N2148,N2162,N2190);
nor #5 GN2149(N2149,N2163,N2193);
nor #5 GN215(N215,N175,N326);
nor #5 GN2150(N2150,N2164,N2196);
nor #5 GN2151(N2151,N2165,N2199);
nor #5 GN2152(N2152,N2166,N2202);
nor #5 GN2153(N2153,N1848,N835);
nor #5 GN2154(N2154,N2031,N662);
nor #5 GN2155(N2155,N1848,N818);
nor #5 GN2156(N2156,N1848,N819);
nor #5 GN2157(N2157,N115,PD5IN);
nor #5 GN2158(N2158,N115,N2157);
nor #5 GN2159(N2159,N2015,N800);
nor #5 GN216(N216,N228,N230);
nor #5 GN2160(N2160,N2017,N801);
nor #5 GN2161(N2161,N2019,N802);
nor #5 GN2162(N2162,N2021,N803);
nor #5 GN2163(N2163,N2023,N804);
nor #5 GN2164(N2164,N2025,N805);
nor #5 GN2165(N2165,N2027,N806);
nor #5 GN2166(N2166,N2029,N807);
nor #5 GN2167(N2167,N1990,N2239);
nor #5 GN2168(N2168,N26,_HD5IN);
nor #5 GN217(N217,N216,N231);
nor #5 GN2172(N2172,N1848,N2157);
nor #5 GN218(N218,N210,N234);
nor #5 GN2181(N2181,N2145,N2272);
nor #5 GN2184(N2184,N2146,N2273);
nor #5 GN2187(N2187,N2147,N2274);
nor #5 GN219(N219,N119,N335);
nor #5 GN2190(N2190,N2148,N2275);
nor #5 GN2193(N2193,N2149,N2276);
nor #5 GN2196(N2196,N2150,N2277);
nor #5 GN2199(N2199,N2151,N2278);
nor #5 GN220(N220,HA2,N39,N40);
nor #5 GN2202(N2202,N2152,N2279);
nor #5 GN221(N221,HA1,N38,N40);
nor #5 GN222(N222,N38,N39,N40);
nor #5 GN223(N223,HA1,HA2,N40);
nor #5 GN2239(N2239,N2168,N26);
nor #5 GN2271(N2271,N2584,N2598);
nor #5 GN2272(N2272,N2159,N800);
nor #5 GN2273(N2273,N2160,N801);
nor #5 GN2274(N2274,N2161,N802);
nor #5 GN2275(N2275,N2162,N803);
nor #5 GN2276(N2276,N2163,N804);
nor #5 GN2277(N2277,N2164,N805);
nor #5 GN2278(N2278,N2165,N806);
nor #5 GN2279(N2279,N2166,N807);
nor #5 GN228(N228,N323,N329,N330);
nor #5 GN2280(N2280,N2271,N601);
nor #5 GN2281(N2281,N2310,N2312);
nor #5 GN2282(N2282,N2281,N510);
nor #5 GN2283(N2283,N2314,N2316);
nor #5 GN2284(N2284,N2283,N579);
nor #5 GN2285(N2285,N2318,N2320);
nor #5 GN2286(N2286,N2285,N581);
nor #5 GN2287(N2287,N2322,N2324);
nor #5 GN2288(N2288,N2287,N583);
nor #5 GN2289(N2289,N2326,N2328);
nor #5 GN2290(N2290,N2289,N585);
nor #5 GN2291(N2291,N2330,N2332);
nor #5 GN2292(N2292,N2291,N587);
nor #5 GN2293(N2293,N2334,N2336);
nor #5 GN2294(N2294,N2293,N589);
nor #5 GN2295(N2295,N2338,N2340);
nor #5 GN2296(N2296,N269,N335);
nor #5 GN2298(N2298,N269,N325);
nor #5 GN2299(N2299,N2438,N2473);
nor #5 GN23(N23,DACK);
nor #5 GN230(N230,N269);
nor #5 GN2300(N2300,N2308,N269);
nor #5 GN2301(N2301,N2295,N498);
nor #5 GN2303(N2303,N2299,N326);
nor #5 GN2306(N2306,N2415,N924);
nor #5 GN2308(N2308,N1206,N2412,N2415);
nor #5 GN231(N231,N256,N269);
nor #5 GN2310(N2310,N2281,N2416);
nor #5 GN2312(N2312,N2570,N701);
nor #5 GN2314(N2314,N2283,N2417);
nor #5 GN2316(N2316,N2571,N702);
nor #5 GN2318(N2318,N2285,N2418);
nor #5 GN2320(N2320,N2572,N703);
nor #5 GN2322(N2322,N2287,N2419);
nor #5 GN2324(N2324,N2573,N704);
nor #5 GN2326(N2326,N2289,N2420);
nor #5 GN2328(N2328,N2574,N705);
nor #5 GN2330(N2330,N2291,N2421);
nor #5 GN2332(N2332,N2575,N706);
nor #5 GN2334(N2334,N2293,N2422);
nor #5 GN2336(N2336,N2576,N707);
nor #5 GN2338(N2338,N2295,N2423);
nor #5 GN234(N234,N269,N320);
nor #5 GN2340(N2340,N2423,N792);
nor #5 GN235(N235,N269);
nor #5 GN237(N237,N333,N347,N436);
nor #5 GN2379(N2379,N2437,N2471);
nor #5 GN2380(N2380,N2457,N2496);
nor #5 GN24(N24,N23,N33,PA0,PA1);
nor #5 GN2412(N2412,N1206,N924);
nor #5 GN2414(N2414,N2379,N327);
nor #5 GN2415(N2415,N2593,N2594);
nor #5 GN2416(N2416,N2312,N701);
nor #5 GN2417(N2417,N2316,N702);
nor #5 GN2418(N2418,N2320,N703);
nor #5 GN2419(N2419,N2324,N704);
nor #5 GN2420(N2420,N2328,N705);
nor #5 GN2421(N2421,N2332,N706);
nor #5 GN2422(N2422,N2336,N707);
nor #5 GN2423(N2423,N2577,N792);
nor #5 GN2424(N2424,N2280,N601);
nor #5 GN2425(N2425,N2282,N510);
nor #5 GN2426(N2426,N2284,N579);
nor #5 GN2427(N2427,N2286,N581);
nor #5 GN2428(N2428,N2288,N583);
nor #5 GN2429(N2429,N2290,N585);
nor #5 GN2430(N2430,N2292,N587);
nor #5 GN2431(N2431,N2294,N589);
nor #5 GN2432(N2432,N2380,N441);
nor #5 GN2433(N2433,N2435,N442);
nor #5 GN2434(N2434,N2436,N2469);
nor #5 GN2435(N2435,N2461,N2565);
nor #5 GN2436(N2436,N2434,N2566);
nor #5 GN2437(N2437,N2379,N2567);
nor #5 GN2438(N2438,N2299,N2568);
nor #5 GN2439(N2439,N2462,N2569);
nor #5 GN2440(N2440,N2280,N2441);
nor #5 GN2441(N2441,N2424,N2440);
nor #5 GN2442(N2442,N2282,N2443);
nor #5 GN2443(N2443,N2425,N2442);
nor #5 GN2444(N2444,N2284,N2445);
nor #5 GN2445(N2445,N2426,N2444);
nor #5 GN2446(N2446,N2286,N2447);
nor #5 GN2447(N2447,N2427,N2446);
nor #5 GN2448(N2448,N2288,N2449);
nor #5 GN2449(N2449,N2428,N2448);
nor #5 GN2450(N2450,N2290,N2451);
nor #5 GN2451(N2451,N2429,N2450);
nor #5 GN2452(N2452,N2292,N2453);
nor #5 GN2453(N2453,N2430,N2452);
nor #5 GN2454(N2454,N2294,N2455);
nor #5 GN2455(N2455,N2431,N2454);
nor #5 GN2456(N2456,N2463,N2578);
nor #5 GN2457(N2457,N2380,N2579);
nor #5 GN2458(N2458,N2459,N2498);
nor #5 GN2459(N2459,N2458,N2580);
nor #5 GN2460(N2460,N2500,N2502);
nor #5 GN2461(N2461,N2435,N2467);
nor #5 GN2462(N2462,N2439,N2475);
nor #5 GN2463(N2463,N2456,N2494);
nor #5 GN2464(N2464,N2458,N496);
nor #5 GN2465(N2465,N2434,N459);
nor #5 GN2467(N2467,N2415,N824);
nor #5 GN2469(N2469,N2566,N808);
nor #5 GN2471(N2471,N2567,N809);
nor #5 GN2473(N2473,N2568,N632);
nor #5 GN2475(N2475,N2569,N338);
nor #5 GN2494(N2494,N2578,N835);
nor #5 GN2496(N2496,N2579,N662);
nor #5 GN2498(N2498,N2580,N818);
nor #5 GN25(N25,N23,N32,N33,PA0);
nor #5 GN2500(N2500,N2460,N2581);
nor #5 GN2502(N2502,N2581,N819);
nor #5 GN2504(N2504,N2460,N334);
nor #5 GN256(N256,N330);
nor #5 GN2565(N2565,N2467,N824);
nor #5 GN2566(N2566,N2415,N808);
nor #5 GN2567(N2567,N2415,N809);
nor #5 GN2568(N2568,N2439,N632);
nor #5 GN2569(N2569,N2415,N338);
nor #5 GN2570(N2570,N2585,N2607);
nor #5 GN2571(N2571,N2586,N2610);
nor #5 GN2572(N2572,N2587,N2613);
nor #5 GN2573(N2573,N2588,N2616);
nor #5 GN2574(N2574,N2589,N2619);
nor #5 GN2575(N2575,N2590,N2622);
nor #5 GN2576(N2576,N2591,N2625);
nor #5 GN2577(N2577,N2592,N2628);
nor #5 GN2578(N2578,N2271,N835);
nor #5 GN2579(N2579,N2456,N662);
nor #5 GN2580(N2580,N2271,N818);
nor #5 GN2581(N2581,N2271,N819);
nor #5 GN2583(N2583,N115,PD4IN);
nor #5 GN2584(N2584,N115,N2583);
nor #5 GN2585(N2585,N2440,N800);
nor #5 GN2586(N2586,N2442,N801);
nor #5 GN2587(N2587,N2444,N802);
nor #5 GN2588(N2588,N2446,N803);
nor #5 GN2589(N2589,N2448,N804);
nor #5 GN2590(N2590,N2450,N805);
nor #5 GN2591(N2591,N2452,N806);
nor #5 GN2592(N2592,N2454,N807);
nor #5 GN2593(N2593,N2415,N2665);
nor #5 GN2594(N2594,N26,_HD4IN);
nor #5 GN2598(N2598,N2271,N2583);
nor #5 GN26(N26,N36);
nor #5 GN2607(N2607,N2570,N2697);
nor #5 GN2610(N2610,N2571,N2698);
nor #5 GN2613(N2613,N2572,N2699);
nor #5 GN2616(N2616,N2573,N2700);
nor #5 GN2619(N2619,N2574,N2701);
nor #5 GN2622(N2622,N2575,N2702);
nor #5 GN2625(N2625,N2576,N2703);
nor #5 GN2628(N2628,N2577,N2704);
nor #5 GN265(N265,N318,N434);
nor #5 GN2665(N2665,N2594,N26);
nor #5 GN269(N269,N2300,N2306,N2412);
nor #5 GN2696(N2696,N2707,N2729);
nor #5 GN2697(N2697,N2585,N800);
nor #5 GN2698(N2698,N2586,N801);
nor #5 GN2699(N2699,N2587,N802);
nor #5 GN27(N27,HA0,N38,N39);
nor #5 GN2700(N2700,N2588,N803);
nor #5 GN2701(N2701,N2589,N804);
nor #5 GN2702(N2702,N2590,N805);
nor #5 GN2703(N2703,N2591,N806);
nor #5 GN2704(N2704,N2592,N807);
nor #5 GN2705(N2705,N2764,N2766);
nor #5 GN2706(N2706,N115,PD3IN);
nor #5 GN2707(N2707,N115,N2706);
nor #5 GN2708(N2708,N2696,N601);
nor #5 GN2709(N2709,N2736,N2738);
nor #5 GN2710(N2710,N2709,N510);
nor #5 GN2711(N2711,N2740,N2742);
nor #5 GN2712(N2712,N2711,N579);
nor #5 GN2713(N2713,N2744,N2746);
nor #5 GN2714(N2714,N2713,N581);
nor #5 GN2715(N2715,N2748,N2750);
nor #5 GN2716(N2716,N2715,N583);
nor #5 GN2717(N2717,N2752,N2754);
nor #5 GN2718(N2718,N2717,N585);
nor #5 GN2719(N2719,N2756,N2758);
nor #5 GN2720(N2720,N2719,N587);
nor #5 GN2721(N2721,N2760,N2762);
nor #5 GN2722(N2722,N2721,N589);
nor #5 GN2723(N2723,N2885,N2927);
nor #5 GN2724(N2724,N1434,N2734);
nor #5 GN2725(N2725,N2723,N496);
nor #5 GN2726(N2726,N2705,N498);
nor #5 GN2729(N2729,N2696,N2706);
nor #5 GN2732(N2732,N2838,N924);
nor #5 GN2734(N2734,N1206,N2837,N2838);
nor #5 GN2736(N2736,N2709,N2839);
nor #5 GN2738(N2738,N2999,N701);
nor #5 GN2740(N2740,N2711,N2840);
nor #5 GN2742(N2742,N3000,N702);
nor #5 GN2744(N2744,N2713,N2841);
nor #5 GN2746(N2746,N3001,N703);
nor #5 GN2748(N2748,N2715,N2842);
nor #5 GN2750(N2750,N3002,N704);
nor #5 GN2752(N2752,N2717,N2843);
nor #5 GN2754(N2754,N3003,N705);
nor #5 GN2756(N2756,N2719,N2844);
nor #5 GN2758(N2758,N3004,N706);
nor #5 GN2760(N2760,N2721,N2845);
nor #5 GN2762(N2762,N3005,N707);
nor #5 GN2764(N2764,N2705,N2846);
nor #5 GN2766(N2766,N2846,N792);
nor #5 GN28(N28,HA0,HA1,N38);
nor #5 GN2837(N2837,N1206,N924);
nor #5 GN2838(N2838,N3020,N3021);
nor #5 GN2839(N2839,N2738,N701);
nor #5 GN2840(N2840,N2742,N702);
nor #5 GN2841(N2841,N2746,N703);
nor #5 GN2842(N2842,N2750,N704);
nor #5 GN2843(N2843,N2754,N705);
nor #5 GN2844(N2844,N2758,N706);
nor #5 GN2845(N2845,N2762,N707);
nor #5 GN2846(N2846,N3006,N792);
nor #5 GN2847(N2847,N2929,N2931);
nor #5 GN2848(N2848,N2708,N601);
nor #5 GN2849(N2849,N2710,N510);
nor #5 GN285(N285,N175,N442);
nor #5 GN2850(N2850,N2712,N579);
nor #5 GN2851(N2851,N2714,N581);
nor #5 GN2852(N2852,N2716,N583);
nor #5 GN2853(N2853,N2718,N585);
nor #5 GN2854(N2854,N2720,N587);
nor #5 GN2855(N2855,N2722,N589);
nor #5 GN2856(N2856,N2847,N334);
nor #5 GN2857(N2857,N1434,N335);
nor #5 GN2859(N2859,N2864,N2902);
nor #5 GN286(N286,N119,N334);
nor #5 GN2861(N2861,N2888,N2994);
nor #5 GN2862(N2862,N2889,N2995);
nor #5 GN2863(N2863,N2890,N2996);
nor #5 GN2864(N2864,N2859,N2997);
nor #5 GN2865(N2865,N2891,N2998);
nor #5 GN2866(N2866,N2708,N2867);
nor #5 GN2867(N2867,N2848,N2866);
nor #5 GN2868(N2868,N2710,N2869);
nor #5 GN2869(N2869,N2849,N2868);
nor #5 GN287(N287,N119,N441);
nor #5 GN2870(N2870,N2712,N2871);
nor #5 GN2871(N2871,N2850,N2870);
nor #5 GN2872(N2872,N2714,N2873);
nor #5 GN2873(N2873,N2851,N2872);
nor #5 GN2874(N2874,N2716,N2875);
nor #5 GN2875(N2875,N2852,N2874);
nor #5 GN2876(N2876,N2718,N2877);
nor #5 GN2877(N2877,N2853,N2876);
nor #5 GN2878(N2878,N2720,N2879);
nor #5 GN2879(N2879,N2854,N2878);
nor #5 GN2880(N2880,N2722,N2881);
nor #5 GN2881(N2881,N2855,N2880);
nor #5 GN2882(N2882,N2892,N3007);
nor #5 GN2883(N2883,N2884,N2925);
nor #5 GN2884(N2884,N2883,N3008);
nor #5 GN2885(N2885,N2723,N3009);
nor #5 GN2887(N2887,N1434,N325);
nor #5 GN2888(N2888,N2861,N2896);
nor #5 GN2889(N2889,N2862,N2898);
nor #5 GN2890(N2890,N2863,N2900);
nor #5 GN2891(N2891,N2865,N2904);
nor #5 GN2892(N2892,N2882,N2923);
nor #5 GN2894(N2894,N2859,N326);
nor #5 GN2896(N2896,N2838,N824);
nor #5 GN2898(N2898,N2995,N808);
nor #5 GN2900(N2900,N2996,N809);
nor #5 GN2902(N2902,N2997,N632);
nor #5 GN2904(N2904,N2998,N338);
nor #5 GN2923(N2923,N3007,N835);
nor #5 GN2925(N2925,N3008,N662);
nor #5 GN2927(N2927,N3009,N818);
nor #5 GN2929(N2929,N2847,N3010);
nor #5 GN2931(N2931,N3010,N819);
nor #5 GN2933(N2933,N2883,N441);
nor #5 GN2993(N2993,N2890,N327);
nor #5 GN2994(N2994,N2896,N824);
nor #5 GN2995(N2995,N2838,N808);
nor #5 GN2996(N2996,N2838,N809);
nor #5 GN2997(N2997,N2865,N632);
nor #5 GN2998(N2998,N2838,N338);
nor #5 GN2999(N2999,N3012,N3033);
nor #5 GN3000(N3000,N3013,N3036);
nor #5 GN3001(N3001,N3014,N3039);
nor #5 GN3002(N3002,N3015,N3042);
nor #5 GN3003(N3003,N3016,N3045);
nor #5 GN3004(N3004,N3017,N3048);
nor #5 GN3005(N3005,N3018,N3051);
nor #5 GN3006(N3006,N3019,N3054);
nor #5 GN3007(N3007,N2696,N835);
nor #5 GN3008(N3008,N2882,N662);
nor #5 GN3009(N3009,N2696,N818);
nor #5 GN3010(N3010,N2696,N819);
nor #5 GN3011(N3011,N2861,N442);
nor #5 GN3012(N3012,N2866,N800);
nor #5 GN3013(N3013,N2868,N801);
nor #5 GN3014(N3014,N2870,N802);
nor #5 GN3015(N3015,N2872,N803);
nor #5 GN3016(N3016,N2874,N804);
nor #5 GN3017(N3017,N2876,N805);
nor #5 GN3018(N3018,N2878,N806);
nor #5 GN3019(N3019,N2880,N807);
nor #5 GN3020(N3020,N2838,N3093);
nor #5 GN3021(N3021,N26,_HD3IN);
nor #5 GN3023(N3023,N2889,N459);
nor #5 GN3033(N3033,N2999,N3125);
nor #5 GN3036(N3036,N3000,N3126);
nor #5 GN3039(N3039,N3001,N3127);
nor #5 GN3042(N3042,N3002,N3128);
nor #5 GN3045(N3045,N3003,N3129);
nor #5 GN3048(N3048,N3004,N3130);
nor #5 GN3051(N3051,N3005,N3131);
nor #5 GN3054(N3054,N3006,N3132);
nor #5 GN3093(N3093,N26,N3021);
nor #5 GN31(N31,PA0);
nor #5 GN3124(N3124,N3441,N3455);
nor #5 GN3125(N3125,N3012,N800);
nor #5 GN3126(N3126,N3013,N801);
nor #5 GN3127(N3127,N3014,N802);
nor #5 GN3128(N3128,N3015,N803);
nor #5 GN3129(N3129,N3016,N804);
nor #5 GN3130(N3130,N3017,N805);
nor #5 GN3131(N3131,N3018,N806);
nor #5 GN3132(N3132,N3019,N807);
nor #5 GN3133(N3133,N3157,N3166,N3270);
nor #5 GN3134(N3134,N1327,N3590);
nor #5 GN3135(N3135,N3124,N601);
nor #5 GN3136(N3136,N3170,N3172);
nor #5 GN3137(N3137,N3136,N510);
nor #5 GN3138(N3138,N3174,N3176);
nor #5 GN3139(N3139,N3138,N579);
nor #5 GN3140(N3140,N3178,N3180);
nor #5 GN3141(N3141,N3140,N581);
nor #5 GN3142(N3142,N3182,N3184);
nor #5 GN3143(N3143,N3142,N583);
nor #5 GN3144(N3144,N3186,N3188);
nor #5 GN3145(N3145,N3144,N585);
nor #5 GN3146(N3146,N3190,N3192);
nor #5 GN3147(N3147,N3146,N587);
nor #5 GN3148(N3148,N3194,N3196);
nor #5 GN3149(N3149,N3148,N589);
nor #5 GN3150(N3150,N3198,N3200);
nor #5 GN3151(N3151,N3133,N335);
nor #5 GN3153(N3153,N3133,N325);
nor #5 GN3154(N3154,N3296,N3331);
nor #5 GN3156(N3156,N1453,N3164);
nor #5 GN3157(N3157,N3133,N3168);
nor #5 GN3158(N3158,N3150,N498);
nor #5 GN3160(N3160,N3154,N326);
nor #5 GN3164(N3164,N3133);
nor #5 GN3166(N3166,N3272,N924);
nor #5 GN3168(N3168,N1206,N3270,N3272);
nor #5 GN317(N317,N372);
nor #5 GN3170(N3170,N3136,N3273);
nor #5 GN3172(N3172,N3428,N701);
nor #5 GN3174(N3174,N3138,N3274);
nor #5 GN3176(N3176,N3429,N702);
nor #5 GN3178(N3178,N3140,N3275);
nor #5 GN318(N318,N217,N265);
nor #5 GN3180(N3180,N3430,N703);
nor #5 GN3182(N3182,N3142,N3276);
nor #5 GN3184(N3184,N3431,N704);
nor #5 GN3186(N3186,N3144,N3277);
nor #5 GN3188(N3188,N3432,N705);
nor #5 GN319(N319,N218,N317,N343);
nor #5 GN3190(N3190,N3146,N3278);
nor #5 GN3192(N3192,N3433,N706);
nor #5 GN3194(N3194,N3148,N3279);
nor #5 GN3196(N3196,N3434,N707);
nor #5 GN3198(N3198,N3150,N3280);
nor #5 GN32(N32,PA1);
nor #5 GN320(N320,N333);
nor #5 GN3200(N3200,N3280,N792);
nor #5 GN321(N321,N265,N319);
nor #5 GN322(N322,N125,N326);
nor #5 GN323(N323,N464,N594);
nor #5 GN3237(N3237,N3295,N3329);
nor #5 GN3238(N3238,N3315,N3354);
nor #5 GN324(N324,N127,N317,N498);
nor #5 GN325(N325,N140);
nor #5 GN326(N326,N213,N23);
nor #5 GN327(N327,N214);
nor #5 GN3270(N3270,N1206,N924);
nor #5 GN3271(N3271,N3237,N327);
nor #5 GN3272(N3272,N3450,N3451);
nor #5 GN3273(N3273,N3172,N701);
nor #5 GN3274(N3274,N3176,N702);
nor #5 GN3275(N3275,N3180,N703);
nor #5 GN3276(N3276,N3184,N704);
nor #5 GN3277(N3277,N3188,N705);
nor #5 GN3278(N3278,N3192,N706);
nor #5 GN3279(N3279,N3196,N707);
nor #5 GN328(N328,N338);
nor #5 GN3280(N3280,N3435,N792);
nor #5 GN3281(N3281,N3135,N601);
nor #5 GN3282(N3282,N3137,N510);
nor #5 GN3283(N3283,N3139,N579);
nor #5 GN3284(N3284,N3141,N581);
nor #5 GN3285(N3285,N3143,N583);
nor #5 GN3286(N3286,N3145,N585);
nor #5 GN3287(N3287,N3147,N587);
nor #5 GN3288(N3288,N3149,N589);
nor #5 GN3289(N3289,N3238,N441);
nor #5 GN329(N329,N328,N592,N594,N632);
nor #5 GN3291(N3291,N3293,N442);
nor #5 GN3292(N3292,N3294,N3327);
nor #5 GN3293(N3293,N3319,N3423);
nor #5 GN3294(N3294,N3292,N3424);
nor #5 GN3295(N3295,N3237,N3425);
nor #5 GN3296(N3296,N3154,N3426);
nor #5 GN3297(N3297,N3320,N3427);
nor #5 GN3298(N3298,N3135,N3299);
nor #5 GN3299(N3299,N3281,N3298);
nor #5 GN33(N33,PA2);
nor #5 GN330(N330,N329,N737);
nor #5 GN3300(N3300,N3137,N3301);
nor #5 GN3301(N3301,N3282,N3300);
nor #5 GN3302(N3302,N3139,N3303);
nor #5 GN3303(N3303,N3283,N3302);
nor #5 GN3304(N3304,N3141,N3305);
nor #5 GN3305(N3305,N3284,N3304);
nor #5 GN3306(N3306,N3143,N3307);
nor #5 GN3307(N3307,N3285,N3306);
nor #5 GN3308(N3308,N3145,N3309);
nor #5 GN3309(N3309,N3286,N3308);
nor #5 GN331(N331,N323);
nor #5 GN3310(N3310,N3147,N3311);
nor #5 GN3311(N3311,N3287,N3310);
nor #5 GN3312(N3312,N3149,N3313);
nor #5 GN3313(N3313,N3288,N3312);
nor #5 GN3314(N3314,N3321,N3436);
nor #5 GN3315(N3315,N3238,N3437);
nor #5 GN3316(N3316,N3317,N3356);
nor #5 GN3317(N3317,N3316,N3438);
nor #5 GN3318(N3318,N3358,N3360);
nor #5 GN3319(N3319,N3293,N3325);
nor #5 GN332(N332,HRST);
nor #5 GN3320(N3320,N3297,N3333);
nor #5 GN3321(N3321,N3314,N3352);
nor #5 GN3322(N3322,N3316,N496);
nor #5 GN3323(N3323,N3292,N459);
nor #5 GN3325(N3325,N3272,N824);
nor #5 GN3327(N3327,N3424,N808);
nor #5 GN3329(N3329,N3425,N809);
nor #5 GN333(N333,N317,N347,N772);
nor #5 GN3331(N3331,N3426,N632);
nor #5 GN3333(N3333,N338,N3427);
nor #5 GN334(N334,N220);
nor #5 GN335(N335,N141);
nor #5 GN3352(N3352,N3436,N835);
nor #5 GN3354(N3354,N3437,N662);
nor #5 GN3356(N3356,N3438,N818);
nor #5 GN3358(N3358,N3318,N3439);
nor #5 GN3360(N3360,N3439,N819);
nor #5 GN3362(N3362,N3318,N334);
nor #5 GN338(N338,N323);
nor #5 GN34(N34,N25);
nor #5 GN3423(N3423,N3325,N824);
nor #5 GN3424(N3424,N3272,N808);
nor #5 GN3425(N3425,N3272,N809);
nor #5 GN3426(N3426,N3297,N632);
nor #5 GN3427(N3427,N3272,N338);
nor #5 GN3428(N3428,N3442,N3464);
nor #5 GN3429(N3429,N3443,N3467);
nor #5 GN343(N343,N319,N398);
nor #5 GN3430(N3430,N3444,N3470);
nor #5 GN3431(N3431,N3445,N3473);
nor #5 GN3432(N3432,N3446,N3476);
nor #5 GN3433(N3433,N3447,N3479);
nor #5 GN3434(N3434,N3448,N3482);
nor #5 GN3435(N3435,N3449,N3485);
nor #5 GN3436(N3436,N3124,N835);
nor #5 GN3437(N3437,N3314,N662);
nor #5 GN3438(N3438,N3124,N818);
nor #5 GN3439(N3439,N3124,N819);
nor #5 GN3440(N3440,N115,PD2IN);
nor #5 GN3441(N3441,N115,N3440);
nor #5 GN3442(N3442,N3298,N800);
nor #5 GN3443(N3443,N3300,N801);
nor #5 GN3444(N3444,N3302,N802);
nor #5 GN3445(N3445,N3304,N803);
nor #5 GN3446(N3446,N3306,N804);
nor #5 GN3447(N3447,N3308,N805);
nor #5 GN3448(N3448,N3310,N806);
nor #5 GN3449(N3449,N3312,N807);
nor #5 GN3450(N3450,N3272,N3522);
nor #5 GN3451(N3451,N26,_HD2IN);
nor #5 GN3455(N3455,N3124,N3440);
nor #5 GN3464(N3464,N3428,N3555);
nor #5 GN3467(N3467,N3429,N3556);
nor #5 GN347(N347,N440,N597,N662,N712);
nor #5 GN3470(N3470,N3430,N3557);
nor #5 GN3473(N3473,N3431,N3558);
nor #5 GN3476(N3476,N3432,N3559);
nor #5 GN3479(N3479,N3433,N3560);
nor #5 GN3482(N3482,N3434,N3561);
nor #5 GN3485(N3485,N3435,N3562);
nor #5 GN35(N35,DACK,PNRDS);
nor #5 GN350(N350,N324,N384,N431);
nor #5 GN3522(N3522,N26,N3451);
nor #5 GN3554(N3554,N3869,N3883);
nor #5 GN3555(N3555,N3442,N800);
nor #5 GN3556(N3556,N3443,N801);
nor #5 GN3557(N3557,N3444,N802);
nor #5 GN3558(N3558,N3445,N803);
nor #5 GN3559(N3559,N3446,N804);
nor #5 GN3560(N3560,N3447,N805);
nor #5 GN3561(N3561,N3448,N806);
nor #5 GN3562(N3562,N3449,N807);
nor #5 GN3563(N3563,N3584,N3592,N3697);
nor #5 GN3564(N3564,N3554,N601);
nor #5 GN3565(N3565,N3596,N3598);
nor #5 GN3566(N3566,N3565,N510);
nor #5 GN3567(N3567,N3600,N3602);
nor #5 GN3568(N3568,N3567,N579);
nor #5 GN3569(N3569,N3604,N3606);
nor #5 GN3570(N3570,N3569,N581);
nor #5 GN3571(N3571,N3608,N3610);
nor #5 GN3572(N3572,N3571,N583);
nor #5 GN3573(N3573,N3612,N3614);
nor #5 GN3574(N3574,N3573,N585);
nor #5 GN3575(N3575,N3616,N3618);
nor #5 GN3576(N3576,N3575,N587);
nor #5 GN3577(N3577,N3620,N3622);
nor #5 GN3578(N3578,N3577,N589);
nor #5 GN3579(N3579,N3624,N3626);
nor #5 GN3580(N3580,N335,N3563);
nor #5 GN3582(N3582,N325,N3563);
nor #5 GN3583(N3583,N3723,N3758);
nor #5 GN3584(N3584,N3563,N3594);
nor #5 GN3585(N3585,N3579,N498);
nor #5 GN3587(N3587,N326,N3583);
nor #5 GN3590(N3590,N3563);
nor #5 GN3592(N3592,N3699,N924);
nor #5 GN3594(N3594,N1206,N3697,N3699);
nor #5 GN3596(N3596,N3565,N3700);
nor #5 GN3598(N3598,N3856,N701);
nor #5 GN36(N36,HCS,HRW,N116);
nor #5 GN3600(N3600,N3567,N3701);
nor #5 GN3602(N3602,N3857,N702);
nor #5 GN3604(N3604,N3569,N3702);
nor #5 GN3606(N3606,N3858,N703);
nor #5 GN3608(N3608,N3571,N3703);
nor #5 GN3610(N3610,N3859,N704);
nor #5 GN3612(N3612,N3573,N3704);
nor #5 GN3614(N3614,N3860,N705);
nor #5 GN3616(N3616,N3575,N3705);
nor #5 GN3618(N3618,N3861,N706);
nor #5 GN3620(N3620,N3577,N3706);
nor #5 GN3622(N3622,N3862,N707);
nor #5 GN3624(N3624,N3579,N3707);
nor #5 GN3626(N3626,N3707,N792);
nor #5 GN364(N364,N454,N507);
nor #5 GN3664(N3664,N3722,N3756);
nor #5 GN3665(N3665,N3742,N3781);
nor #5 GN3697(N3697,N1206,N924);
nor #5 GN3698(N3698,N327,N3664);
nor #5 GN3699(N3699,N3878,N3879);
nor #5 GN37(N37,N27);
nor #5 GN3700(N3700,N3598,N701);
nor #5 GN3701(N3701,N3602,N702);
nor #5 GN3702(N3702,N3606,N703);
nor #5 GN3703(N3703,N3610,N704);
nor #5 GN3704(N3704,N3614,N705);
nor #5 GN3705(N3705,N3618,N706);
nor #5 GN3706(N3706,N3622,N707);
nor #5 GN3707(N3707,N3863,N792);
nor #5 GN3708(N3708,N3564,N601);
nor #5 GN3709(N3709,N3566,N510);
nor #5 GN3710(N3710,N3568,N579);
nor #5 GN3711(N3711,N3570,N581);
nor #5 GN3712(N3712,N3572,N583);
nor #5 GN3713(N3713,N3574,N585);
nor #5 GN3714(N3714,N3576,N587);
nor #5 GN3715(N3715,N3578,N589);
nor #5 GN3716(N3716,N3665,N441);
nor #5 GN3718(N3718,N3720,N442);
nor #5 GN3719(N3719,N3721,N3754);
nor #5 GN372(N372,N332,N435);
nor #5 GN3720(N3720,N3746,N3851);
nor #5 GN3721(N3721,N3719,N3852);
nor #5 GN3722(N3722,N3664,N3853);
nor #5 GN3723(N3723,N3583,N3854);
nor #5 GN3724(N3724,N3747,N3855);
nor #5 GN3725(N3725,N3564,N3726);
nor #5 GN3726(N3726,N3708,N3725);
nor #5 GN3727(N3727,N3566,N3728);
nor #5 GN3728(N3728,N3709,N3727);
nor #5 GN3729(N3729,N3568,N3730);
nor #5 GN3730(N3730,N3710,N3729);
nor #5 GN3731(N3731,N3570,N3732);
nor #5 GN3732(N3732,N3711,N3731);
nor #5 GN3733(N3733,N3572,N3734);
nor #5 GN3734(N3734,N3712,N3733);
nor #5 GN3735(N3735,N3574,N3736);
nor #5 GN3736(N3736,N3713,N3735);
nor #5 GN3737(N3737,N3576,N3738);
nor #5 GN3738(N3738,N3714,N3737);
nor #5 GN3739(N3739,N3578,N3740);
nor #5 GN3740(N3740,N3715,N3739);
nor #5 GN3741(N3741,N3748,N3864);
nor #5 GN3742(N3742,N3665,N3865);
nor #5 GN3743(N3743,N3744,N3783);
nor #5 GN3744(N3744,N3743,N3866);
nor #5 GN3745(N3745,N3785,N3787);
nor #5 GN3746(N3746,N3720,N3752);
nor #5 GN3747(N3747,N3724,N3760);
nor #5 GN3748(N3748,N3741,N3779);
nor #5 GN3749(N3749,N3743,N496);
nor #5 GN3750(N3750,N3719,N459);
nor #5 GN3752(N3752,N3699,N824);
nor #5 GN3754(N3754,N3852,N808);
nor #5 GN3756(N3756,N3853,N809);
nor #5 GN3758(N3758,N3854,N632);
nor #5 GN3760(N3760,N338,N3855);
nor #5 GN3779(N3779,N3864,N835);
nor #5 GN3781(N3781,N3865,N662);
nor #5 GN3783(N3783,N3866,N818);
nor #5 GN3785(N3785,N3745,N3867);
nor #5 GN3787(N3787,N3867,N819);
nor #5 GN3789(N3789,N334,N3745);
nor #5 GN38(N38,HA2);
nor #5 GN384(N384,N350,N437);
nor #5 GN3851(N3851,N3752,N824);
nor #5 GN3852(N3852,N3699,N808);
nor #5 GN3853(N3853,N3699,N809);
nor #5 GN3854(N3854,N3724,N632);
nor #5 GN3855(N3855,N338,N3699);
nor #5 GN3856(N3856,N3870,N3892);
nor #5 GN3857(N3857,N3871,N3895);
nor #5 GN3858(N3858,N3872,N3898);
nor #5 GN3859(N3859,N3873,N3901);
nor #5 GN3860(N3860,N3874,N3904);
nor #5 GN3861(N3861,N3875,N3907);
nor #5 GN3862(N3862,N3876,N3910);
nor #5 GN3863(N3863,N3877,N3913);
nor #5 GN3864(N3864,N3554,N835);
nor #5 GN3865(N3865,N3741,N662);
nor #5 GN3866(N3866,N3554,N818);
nor #5 GN3867(N3867,N3554,N819);
nor #5 GN3868(N3868,N115,PD1IN);
nor #5 GN3869(N3869,N115,N3868);
nor #5 GN3870(N3870,N3725,N800);
nor #5 GN3871(N3871,N3727,N801);
nor #5 GN3872(N3872,N3729,N802);
nor #5 GN3873(N3873,N3731,N803);
nor #5 GN3874(N3874,N3733,N804);
nor #5 GN3875(N3875,N3735,N805);
nor #5 GN3876(N3876,N3737,N806);
nor #5 GN3877(N3877,N3739,N807);
nor #5 GN3878(N3878,N3699,N3950);
nor #5 GN3879(N3879,N26,_HD1IN);
nor #5 GN3883(N3883,N3554,N3868);
nor #5 GN3892(N3892,N3856,N3983);
nor #5 GN3895(N3895,N3857,N3984);
nor #5 GN3898(N3898,N3858,N3985);
nor #5 GN39(N39,HA1);
nor #5 GN390(N390,N438,N493);
nor #5 GN3901(N3901,N3859,N3986);
nor #5 GN3904(N3904,N3860,N3987);
nor #5 GN3907(N3907,N3861,N3988);
nor #5 GN3910(N3910,N3862,N3989);
nor #5 GN3913(N3913,N3863,N3990);
nor #5 GN3950(N3950,N26,N3879);
nor #5 GN397(N397,N364,N433);
nor #5 GN398(N398,N320,N399);
nor #5 GN3982(N3982,N4304,N4307);
nor #5 GN3983(N3983,N3870,N800);
nor #5 GN3984(N3984,N3871,N801);
nor #5 GN3985(N3985,N3872,N802);
nor #5 GN3986(N3986,N3873,N803);
nor #5 GN3987(N3987,N3874,N804);
nor #5 GN3988(N3988,N3875,N805);
nor #5 GN3989(N3989,N3876,N806);
nor #5 GN399(N399,N436);
nor #5 GN3990(N3990,N3877,N807);
nor #5 GN3991(N3991,N3982,N601);
nor #5 GN3992(N3992,N4021,N4023);
nor #5 GN3993(N3993,N3992,N510);
nor #5 GN3994(N3994,N4025,N4027);
nor #5 GN3995(N3995,N3994,N579);
nor #5 GN3996(N3996,N4029,N4031);
nor #5 GN3997(N3997,N3996,N581);
nor #5 GN3998(N3998,N4033,N4035);
nor #5 GN3999(N3999,N3998,N583);
nor #5 GN40(N40,HA0);
nor #5 GN4000(N4000,N4037,N4039);
nor #5 GN4001(N4001,N4000,N585);
nor #5 GN4002(N4002,N4041,N4043);
nor #5 GN4003(N4003,N4002,N587);
nor #5 GN4004(N4004,N4045,N4047);
nor #5 GN4005(N4005,N4004,N589);
nor #5 GN4006(N4006,N4049,N4051);
nor #5 GN4007(N4007,N1346,N335);
nor #5 GN4009(N4009,N1346,N325);
nor #5 GN4010(N4010,N4149,N4184);
nor #5 GN4011(N4011,N1346,N4019);
nor #5 GN4012(N4012,N4006,N498);
nor #5 GN4014(N4014,N326,N4010);
nor #5 GN4017(N4017,N4125,N924);
nor #5 GN4019(N4019,N1206,N4123,N4125);
nor #5 GN4021(N4021,N3992,N4126);
nor #5 GN4023(N4023,N4281,N701);
nor #5 GN4025(N4025,N3994,N4127);
nor #5 GN4027(N4027,N4282,N702);
nor #5 GN4029(N4029,N3996,N4128);
nor #5 GN4031(N4031,N4283,N703);
nor #5 GN4033(N4033,N3998,N4129);
nor #5 GN4035(N4035,N4284,N704);
nor #5 GN4037(N4037,N4000,N4130);
nor #5 GN4039(N4039,N4285,N705);
nor #5 GN4041(N4041,N4002,N4131);
nor #5 GN4043(N4043,N4286,N706);
nor #5 GN4045(N4045,N4004,N4132);
nor #5 GN4047(N4047,N4287,N707);
nor #5 GN4049(N4049,N4006,N4133);
nor #5 GN4051(N4051,N4133,N792);
nor #5 GN4090(N4090,N4148,N4182);
nor #5 GN4091(N4091,N4168,N4207);
nor #5 GN4123(N4123,N1206,N924);
nor #5 GN4124(N4124,N327,N4090);
nor #5 GN4125(N4125,N4302,N4303);
nor #5 GN4126(N4126,N4023,N701);
nor #5 GN4127(N4127,N4027,N702);
nor #5 GN4128(N4128,N4031,N703);
nor #5 GN4129(N4129,N4035,N704);
nor #5 GN4130(N4130,N4039,N705);
nor #5 GN4131(N4131,N4043,N706);
nor #5 GN4132(N4132,N4047,N707);
nor #5 GN4133(N4133,N4288,N792);
nor #5 GN4134(N4134,N3991,N601);
nor #5 GN4135(N4135,N3993,N510);
nor #5 GN4136(N4136,N3995,N579);
nor #5 GN4137(N4137,N3997,N581);
nor #5 GN4138(N4138,N3999,N583);
nor #5 GN4139(N4139,N4001,N585);
nor #5 GN4140(N4140,N4003,N587);
nor #5 GN4141(N4141,N4005,N589);
nor #5 GN4142(N4142,N4091,N441);
nor #5 GN4144(N4144,N4146,N442);
nor #5 GN4145(N4145,N4147,N4180);
nor #5 GN4146(N4146,N4172,N4276);
nor #5 GN4147(N4147,N4145,N4277);
nor #5 GN4148(N4148,N4090,N4278);
nor #5 GN4149(N4149,N4010,N4279);
nor #5 GN4150(N4150,N4173,N4280);
nor #5 GN4151(N4151,N3991,N4152);
nor #5 GN4152(N4152,N4134,N4151);
nor #5 GN4153(N4153,N3993,N4154);
nor #5 GN4154(N4154,N4135,N4153);
nor #5 GN4155(N4155,N3995,N4156);
nor #5 GN4156(N4156,N4136,N4155);
nor #5 GN4157(N4157,N3997,N4158);
nor #5 GN4158(N4158,N4137,N4157);
nor #5 GN4159(N4159,N3999,N4160);
nor #5 GN4160(N4160,N4138,N4159);
nor #5 GN4161(N4161,N4001,N4162);
nor #5 GN4162(N4162,N4139,N4161);
nor #5 GN4163(N4163,N4003,N4164);
nor #5 GN4164(N4164,N4140,N4163);
nor #5 GN4165(N4165,N4005,N4166);
nor #5 GN4166(N4166,N4141,N4165);
nor #5 GN4167(N4167,N4174,N4289);
nor #5 GN4168(N4168,N4091,N4290);
nor #5 GN4169(N4169,N4170,N4209);
nor #5 GN4170(N4170,N4169,N4291);
nor #5 GN4171(N4171,N4211,N4213);
nor #5 GN4172(N4172,N4146,N4178);
nor #5 GN4173(N4173,N4150,N4186);
nor #5 GN4174(N4174,N4167,N4205);
nor #5 GN4175(N4175,N4169,N496);
nor #5 GN4176(N4176,N4145,N459);
nor #5 GN4178(N4178,N4125,N824);
nor #5 GN4180(N4180,N4277,N808);
nor #5 GN4182(N4182,N4278,N809);
nor #5 GN4184(N4184,N4279,N632);
nor #5 GN4186(N4186,N338,N4280);
nor #5 GN4205(N4205,N4289,N835);
nor #5 GN4207(N4207,N4290,N662);
nor #5 GN4209(N4209,N4291,N818);
nor #5 GN4211(N4211,N4171,N4292);
nor #5 GN4213(N4213,N4292,N819);
nor #5 GN4215(N4215,N334,N4171);
nor #5 GN4276(N4276,N4178,N824);
nor #5 GN4277(N4277,N4125,N808);
nor #5 GN4278(N4278,N4125,N809);
nor #5 GN4279(N4279,N4150,N632);
nor #5 GN4280(N4280,N338,N4125);
nor #5 GN4281(N4281,N4294,N4316);
nor #5 GN4282(N4282,N4295,N4319);
nor #5 GN4283(N4283,N4296,N4322);
nor #5 GN4284(N4284,N4297,N4325);
nor #5 GN4285(N4285,N4298,N4328);
nor #5 GN4286(N4286,N4299,N4331);
nor #5 GN4287(N4287,N4300,N4334);
nor #5 GN4288(N4288,N4301,N4337);
nor #5 GN4289(N4289,N3982,N835);
nor #5 GN4290(N4290,N4167,N662);
nor #5 GN4291(N4291,N3982,N818);
nor #5 GN4292(N4292,N3982,N819);
nor #5 GN4293(N4293,N115,PD0IN);
nor #5 GN4294(N4294,N4151,N800);
nor #5 GN4295(N4295,N4153,N801);
nor #5 GN4296(N4296,N4155,N802);
nor #5 GN4297(N4297,N4157,N803);
nor #5 GN4298(N4298,N4159,N804);
nor #5 GN4299(N4299,N4161,N805);
nor #5 GN430(N430,N317);
nor #5 GN4300(N4300,N4163,N806);
nor #5 GN4301(N4301,N4165,N807);
nor #5 GN4302(N4302,N26,_HD0IN);
nor #5 GN4303(N4303,N4125,N4375);
nor #5 GN4304(N4304,N115,N4293);
nor #5 GN4307(N4307,N3982,N4293);
nor #5 GN431(N431,N116,N430);
nor #5 GN4316(N4316,N4281,N4406);
nor #5 GN4319(N4319,N4282,N4407);
nor #5 GN432(N432,N322,N439);
nor #5 GN4322(N4322,N4283,N4408);
nor #5 GN4325(N4325,N4284,N4409);
nor #5 GN4328(N4328,N4285,N4410);
nor #5 GN433(N433,N285,N397);
nor #5 GN4331(N4331,N4286,N4411);
nor #5 GN4334(N4334,N4287,N4412);
nor #5 GN4337(N4337,N4288,N4413);
nor #5 GN434(N434,N256,N331);
nor #5 GN435(N435,N1457,N1464,N1570);
nor #5 GN436(N436,N490,N597);
nor #5 GN437(N437,N602,N659);
nor #5 GN4375(N4375,N26,N4302);
nor #5 GN438(N438,N127,N441);
nor #5 GN439(N439,N330,N432);
nor #5 GN440(N440,N390,N438);
nor #5 GN4406(N4406,N4294,N800);
nor #5 GN4407(N4407,N4295,N801);
nor #5 GN4408(N4408,N4296,N802);
nor #5 GN4409(N4409,N4297,N803);
nor #5 GN441(N441,N221);
nor #5 GN4410(N4410,N4298,N804);
nor #5 GN4411(N4411,N4299,N805);
nor #5 GN4412(N4412,N4300,N806);
nor #5 GN4413(N4413,N4301,N807);
nor #5 GN442(N442,N211);
nor #5 GN443(N443,N462,N464);
nor #5 GN444(N444,N285,N433,N507);
nor #5 GN445(N445,N455,N468,N510,N591);
nor #5 GN446(N446,N470,N472,N514,N579);
nor #5 GN447(N447,N473,N475,N518,N581);
nor #5 GN448(N448,N476,N478,N522,N583);
nor #5 GN449(N449,N479,N481,N526,N585);
nor #5 GN450(N450,N456,N483,N530,N587);
nor #5 GN451(N451,N486,N488,N533,N589);
nor #5 GN452(N452,N490,N492);
nor #5 GN453(N453,N219,N466);
nor #5 GN454(N454,N364,N444);
nor #5 GN455(N455,N445,N507,N638,N701);
nor #5 GN456(N456,N450,N526,N653,N706);
nor #5 GN457(N457,N324,N350);
nor #5 GN459(N459,N212);
nor #5 GN462(N462,N287,N443);
nor #5 GN464(N464,N323,N329);
nor #5 GN466(N466,N453,N595,N596);
nor #5 GN468(N468,N455,N717);
nor #5 GN470(N470,N472,N718);
nor #5 GN472(N472,N446,N591,N641,N702);
nor #5 GN473(N473,N475,N719);
nor #5 GN475(N475,N447,N514,N644,N703);
nor #5 GN476(N476,N478,N720);
nor #5 GN478(N478,N448,N518,N647,N704);
nor #5 GN479(N479,N481,N721);
nor #5 GN481(N481,N449,N522,N650,N705);
nor #5 GN483(N483,N456,N722);
nor #5 GN486(N486,N488,N723);
nor #5 GN488(N488,N451,N530,N656,N707);
nor #5 GN490(N490,N317,N347,N436);
nor #5 GN492(N492,N215,N452);
nor #5 GN493(N493,N333,N390);
nor #5 GN496(N496,N222);
nor #5 GN498(N498,N223);
nor #5 GN50(N50,HRW);
nor #5 GN507(N507,N444,N454,N455,N800);
nor #5 GN510(N510,N541);
nor #5 GN514(N514,N446,N475,N542,N802);
nor #5 GN518(N518,N447,N478,N543,N803);
nor #5 GN522(N522,N448,N481,N544,N804);
nor #5 GN526(N526,N449,N456,N545,N805);
nor #5 GN530(N530,N450,N488,N546,N806);
nor #5 GN533(N533,N451,N547,N602,N807);
nor #5 GN541(N541,N445,N578);
nor #5 GN542(N542,N446,N580);
nor #5 GN543(N543,N447,N582);
nor #5 GN544(N544,N448,N584);
nor #5 GN545(N545,N449,N586);
nor #5 GN546(N546,N450,N588);
nor #5 GN547(N547,N451,N590);
nor #5 GN578(N578,N541,N591);
nor #5 GN579(N579,N542);
nor #5 GN580(N580,N514,N542);
nor #5 GN581(N581,N543);
nor #5 GN582(N582,N518,N543);
nor #5 GN583(N583,N544);
nor #5 GN584(N584,N522,N544);
nor #5 GN585(N585,N545);
nor #5 GN586(N586,N526,N545);
nor #5 GN587(N587,N546);
nor #5 GN588(N588,N530,N546);
nor #5 GN589(N589,N547);
nor #5 GN590(N590,N533,N547);
nor #5 GN591(N591,N445,N472,N541,N801);
nor #5 GN592(N592,N322,N432);
nor #5 GN594(N594,N287,N329,N462);
nor #5 GN595(N595,N219,N710,N799);
nor #5 GN596(N596,N219,N716,N799);
nor #5 GN597(N597,N215,N347,N492);
nor #5 GN598(N598,N125,N442);
nor #5 GN599(N599,N125,N459);
nor #5 GN600(N600,N125,N327);
nor #5 GN601(N601,N454);
nor #5 GN602(N602,N457,N533,N659,N711);
nor #5 GN603(N603,N127,N334);
nor #5 GN604(N604,N127,N496);
nor #5 GN628(N628,N317,N599,N714);
nor #5 GN632(N632,N330);
nor #5 GN638(N638,N507,N827);
nor #5 GN641(N641,N591,N828);
nor #5 GN644(N644,N514,N829);
nor #5 GN647(N647,N518,N830);
nor #5 GN650(N650,N522,N831);
nor #5 GN653(N653,N526,N832);
nor #5 GN656(N656,N530,N833);
nor #5 GN659(N659,N437,N457);
nor #5 GN662(N662,N333);
nor #5 GN664(N664,N317,N604,N724);
nor #5 GN666(N666,N317,N603,N725);
nor #5 GN701(N701,N468);
nor #5 GN702(N702,N470);
nor #5 GN703(N703,N473);
nor #5 GN704(N704,N476);
nor #5 GN705(N705,N479);
nor #5 GN706(N706,N483);
nor #5 GN707(N707,N486);
nor #5 GN708(N708,N317,N598,N713);
nor #5 GN709(N709,N317,N600,N715);
nor #5 GN710(N710,N825,N826);
nor #5 GN711(N711,N533,N834);
nor #5 GN712(N712,N835);
nor #5 GN713(N713,N207,N708);
nor #5 GN714(N714,N286,N628);
nor #5 GN715(N715,N208,N709);
nor #5 GN716(N716,N710);
nor #5 GN717(N717,N445,N468);
nor #5 GN718(N718,N446,N470);
nor #5 GN719(N719,N447,N473);
nor #5 GN720(N720,N448,N476);
nor #5 GN721(N721,N449,N479);
nor #5 GN722(N722,N450,N483);
nor #5 GN723(N723,N451,N486);
nor #5 GN724(N724,N209,N664);
nor #5 GN725(N725,N177,N666);
nor #5 GN737(N737,N317,N330,N592);
nor #5 GN772(N772,N333,N440);
nor #5 GN792(N792,N437);
nor #5 GN799(N799,N902);
nor #5 GN800(N800,N638);
nor #5 GN801(N801,N641);
nor #5 GN802(N802,N644);
nor #5 GN803(N803,N647);
nor #5 GN804(N804,N650);
nor #5 GN805(N805,N653);
nor #5 GN806(N806,N656);
nor #5 GN807(N807,N711);
nor #5 GN808(N808,N286);
nor #5 GN809(N809,N208);
nor #5 GN818(N818,N209);
nor #5 GN819(N819,N177);
nor #5 GN822(N822,N115,N837);
nor #5 GN823(N823,N822,N839);
nor #5 GN824(N824,N207);
nor #5 GN825(N825,N710,N876);
nor #5 GN826(N826,N26,_HD7IN);
nor #5 GN827(N827,N455,N638);
nor #5 GN828(N828,N472,N641);
nor #5 GN829(N829,N475,N644);
nor #5 GN830(N830,N478,N647);
nor #5 GN831(N831,N481,N650);
nor #5 GN832(N832,N456,N653);
nor #5 GN833(N833,N488,N656);
nor #5 GN834(N834,N602,N711);
nor #5 GN835(N835,N436);
nor #5 GN837(N837,N115,PD7IN);
nor #5 GN839(N839,N823,N837);
nor #5 GN84(N84,N28);
nor #5 GN876(N876,N26,N826);
nor #5 GN899(N899,N117,N666);
nor #5 GN900(N900,N326,N923);
nor #5 GN901(N901,N974);
nor #5 GN902(N902,N901);
nor #5 GN903(N903,N453);
nor #5 GN904(N904,N601,N823);
nor #5 GN905(N905,N932,N934);
nor #5 GN906(N906,N510,N905);
nor #5 GN907(N907,N936,N938);
nor #5 GN908(N908,N579,N907);
nor #5 GN909(N909,N940,N942);
nor #5 GN910(N910,N581,N909);
nor #5 GN911(N911,N944,N946);
nor #5 GN912(N912,N583,N911);
nor #5 GN913(N913,N948,N950);
nor #5 GN914(N914,N585,N913);
nor #5 GN915(N915,N952,N954);
nor #5 GN916(N916,N587,N915);
nor #5 GN917(N917,N956,N958);
nor #5 GN918(N918,N589,N917);
nor #5 GN919(N919,N960,N962);
nor #5 GN920(N920,N1081,N1119);
nor #5 GN921(N921,N496,N920);
nor #5 GN922(N922,N325,N708);
nor #5 GN923(N923,N1061,N1095);
nor #5 GN924(N924,N332,N596);
nor #5 GN926(N926,N1002,N327);
nor #5 GN932(N932,N1037,N905);
nor #5 GN934(N934,N1194,N701);
nor #5 GN936(N936,N1038,N907);
nor #5 GN938(N938,N1195,N702);
nor #5 GN940(N940,N1039,N909);
nor #5 GN942(N942,N1196,N703);
nor #5 GN944(N944,N1040,N911);
nor #5 GN946(N946,N1197,N704);
nor #5 GN948(N948,N1041,N913);
nor #5 GN950(N950,N1198,N705);
nor #5 GN952(N952,N1042,N915);
nor #5 GN954(N954,N1199,N706);
nor #5 GN956(N956,N1043,N917);
nor #5 GN958(N958,N1200,N707);
nor #5 GN960(N960,N1044,N919);
nor #5 GN962(N962,N1044,N792);
nor #5 GN967(N967,N335,N792);
nor #5 GN974(N974,N1003);
nor #5 GPD0OUT(PD0OUT,N4009,N4014,N4124,N4144,N4176);
nor #5 GPD1OUT(PD1OUT,N3582,N3587,N3698,N3718,N3750);
nor #5 GPD2OUT(PD2OUT,N3153,N3160,N3271,N3291,N3323);
nor #5 GPD3OUT(PD3OUT,N2887,N2894,N2993,N3011,N3023);
nor #5 GPD4OUT(PD4OUT,N2298,N2303,N2414,N2433,N2465);
nor #5 GPD5OUT(PD5OUT,N1874,N1879,N1989,N2008,N2040);
nor #5 GPD6OUT(PD6OUT,N1328,N1329,N1398,N1435,N1455,N1536,N1616,N1688);
nor #5 GPD7OUT(PD7OUT,N1036,N1056,N1087,N1126,N1188,N900,N922,N926);
nor #5 GPDOEA(PDOEA,DACK,PNWDS);
nor #5 GPDOEB(PDOEB,PCS,PNRDS);
nor #5 GPIRQ(PIRQ,N3134,N3156);
nor #5 GPNMI(PNMI,N1332);
nor #5 GPRST(PRST,N1433,N332);
nor #5 inv_HD0IN(_HD0IN,HD0IN);
nor #5 inv_HD1IN(_HD1IN,HD1IN);
nor #5 inv_HD2IN(_HD2IN,HD2IN);
nor #5 inv_HD3IN(_HD3IN,HD3IN);
nor #5 inv_HD4IN(_HD4IN,HD4IN);
nor #5 inv_HD5IN(_HD5IN,HD5IN);
nor #5 inv_HD6IN(_HD6IN,HD6IN);
nor #5 inv_HD7IN(_HD7IN,HD7IN);
nor #5 nor_hdoe(HDOE,HDOEA);
nor #5 nor_pdoe(PDOE,PDOEA,PDOEB);
endmodule
