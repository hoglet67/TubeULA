module tube_ula(
      DACK
    , DRQ
    , HA0
    , HA1
    , HA2
    , HCS
    , HD0IN
    , HD0OUT
    , HD1IN
    , HD1OUT
    , HD2IN
    , HD2OUT
    , HD3IN
    , HD3OUT
    , HD4IN
    , HD4OUT
    , HD5IN
    , HD5OUT
    , HD6IN
    , HD6OUT
    , HD7IN
    , HD7OUT
    , HDOE
    , HDOEA
    , HIRQ
    , HO2
    , HRST
    , HRW
    , PA0
    , PA1
    , PA2
    , PCS
    , PD0IN
    , PD0OUT
    , PD1IN
    , PD1OUT
    , PD2IN
    , PD2OUT
    , PD3IN
    , PD3OUT
    , PD4IN
    , PD4OUT
    , PD5IN
    , PD5OUT
    , PD6IN
    , PD6OUT
    , PD7IN
    , PD7OUT
    , PDOE
    , PDOEA
    , PDOEB
    , PIRQ
    , PNMI
    , PNRDS
    , PNWDS
    , PRST
);
// Inputs
input DACK;
input HA0;
input HA1;
input HA2;
input HCS;
input HD0IN;
input HD1IN;
input HD2IN;
input HD3IN;
input HD4IN;
input HD5IN;
input HD6IN;
input HD7IN;
input HO2;
input HRST;
input HRW;
input PA0;
input PA1;
input PA2;
input PCS;
input PD0IN;
input PD1IN;
input PD2IN;
input PD3IN;
input PD4IN;
input PD5IN;
input PD6IN;
input PD7IN;
input PNRDS;
input PNWDS;
// Outputs
output DRQ;
output HD0OUT;
output HD1OUT;
output HD2OUT;
output HD3OUT;
output HD4OUT;
output HD5OUT;
output HD6OUT;
output HD7OUT;
output HDOE;
output HDOEA;
output HIRQ;
output PD0OUT;
output PD1OUT;
output PD2OUT;
output PD3OUT;
output PD4OUT;
output PD5OUT;
output PD6OUT;
output PD7OUT;
output PDOE;
output PDOEA;
output PDOEB;
output PIRQ;
output PNMI;
output PRST;
// Wires
wire N1002;
wire N1003;
wire N1004;
wire N1035;
wire N1036;
wire N1056;
wire N1057;
wire N1058;
wire N1059;
wire N1060;
wire N1061;
wire N1062;
wire N1063;
wire N1064;
wire N1065;
wire N1066;
wire N1067;
wire N1068;
wire N1069;
wire N1070;
wire N1071;
wire N1072;
wire N1073;
wire N1074;
wire N1075;
wire N1076;
wire N1077;
wire N1078;
wire N1079;
wire N1080;
wire N1081;
wire N1082;
wire N1083;
wire N1084;
wire N1085;
wire N1086;
wire N1087;
wire N1121;
wire N1125;
wire N1126;
wire N115;
wire N1155;
wire N116;
wire N117;
wire N118;
wire N1187;
wire N1188;
wire N119;
wire N1194;
wire N1195;
wire N1196;
wire N1197;
wire N1198;
wire N1199;
wire N120;
wire N1200;
wire N1201;
wire N1206;
wire N1208;
wire N121;
wire N122;
wire N1226;
wire N1229;
wire N123;
wire N1232;
wire N1235;
wire N1238;
wire N124;
wire N1241;
wire N1244;
wire N1247;
wire N125;
wire N126;
wire N127;
wire N1314;
wire N1326;
wire N1327;
wire N1328;
wire N1329;
wire N1332;
wire N1335;
wire N1336;
wire N1339;
wire N1343;
wire N1346;
wire N1349;
wire N1396;
wire N1398;
wire N1399;
wire N140;
wire N141;
wire N1430;
wire N1431;
wire N1432;
wire N1433;
wire N1434;
wire N1435;
wire N1436;
wire N1437;
wire N1439;
wire N1441;
wire N1443;
wire N1445;
wire N1447;
wire N1449;
wire N1451;
wire N1453;
wire N1455;
wire N1456;
wire N1457;
wire N1458;
wire N1464;
wire N1466;
wire N1468;
wire N1472;
wire N1476;
wire N1480;
wire N1484;
wire N1488;
wire N1492;
wire N1496;
wire N1536;
wire N1537;
wire N1538;
wire N1570;
wire N1571;
wire N1588;
wire N1589;
wire N1590;
wire N1591;
wire N1592;
wire N1593;
wire N1594;
wire N1595;
wire N1596;
wire N1597;
wire N1598;
wire N1599;
wire N1600;
wire N1601;
wire N1602;
wire N1603;
wire N1604;
wire N1605;
wire N1606;
wire N1607;
wire N1608;
wire N1609;
wire N1610;
wire N1611;
wire N1612;
wire N1613;
wire N1614;
wire N1616;
wire N1617;
wire N1618;
wire N1619;
wire N1620;
wire N1655;
wire N1687;
wire N1688;
wire N1724;
wire N1725;
wire N1726;
wire N1727;
wire N1728;
wire N1729;
wire N1730;
wire N1731;
wire N1745;
wire N175;
wire N1750;
wire N1759;
wire N176;
wire N1762;
wire N1765;
wire N1768;
wire N177;
wire N1771;
wire N1774;
wire N1777;
wire N1780;
wire N1848;
wire N1858;
wire N1860;
wire N1862;
wire N1864;
wire N1866;
wire N1868;
wire N1870;
wire N1872;
wire N1873;
wire N1874;
wire N1875;
wire N1876;
wire N1877;
wire N1879;
wire N1882;
wire N1884;
wire N1886;
wire N1890;
wire N1894;
wire N1898;
wire N1902;
wire N1906;
wire N1910;
wire N1914;
wire N1955;
wire N1956;
wire N1988;
wire N1989;
wire N1990;
wire N2007;
wire N2008;
wire N2009;
wire N2010;
wire N2011;
wire N2012;
wire N2013;
wire N2014;
wire N2015;
wire N2016;
wire N2017;
wire N2018;
wire N2019;
wire N2020;
wire N2021;
wire N2022;
wire N2023;
wire N2024;
wire N2025;
wire N2026;
wire N2027;
wire N2028;
wire N2029;
wire N2030;
wire N2031;
wire N2032;
wire N2033;
wire N2034;
wire N2035;
wire N2036;
wire N2037;
wire N2038;
wire N2039;
wire N2040;
wire N207;
wire N2075;
wire N2079;
wire N208;
wire N209;
wire N210;
wire N211;
wire N212;
wire N213;
wire N214;
wire N2145;
wire N2146;
wire N2147;
wire N2148;
wire N2149;
wire N215;
wire N2150;
wire N2151;
wire N2152;
wire N216;
wire N2167;
wire N217;
wire N2172;
wire N218;
wire N2181;
wire N2184;
wire N2187;
wire N219;
wire N2190;
wire N2193;
wire N2196;
wire N2199;
wire N220;
wire N2202;
wire N221;
wire N222;
wire N223;
wire N2271;
wire N228;
wire N2281;
wire N2283;
wire N2285;
wire N2287;
wire N2289;
wire N2291;
wire N2293;
wire N2295;
wire N2296;
wire N2298;
wire N2299;
wire N23;
wire N230;
wire N2300;
wire N2301;
wire N2303;
wire N2306;
wire N2308;
wire N231;
wire N2310;
wire N2314;
wire N2318;
wire N2322;
wire N2326;
wire N2330;
wire N2334;
wire N2338;
wire N234;
wire N235;
wire N237;
wire N2379;
wire N2380;
wire N24;
wire N2412;
wire N2414;
wire N2415;
wire N2432;
wire N2433;
wire N2434;
wire N2435;
wire N2436;
wire N2437;
wire N2438;
wire N2439;
wire N2440;
wire N2441;
wire N2442;
wire N2443;
wire N2444;
wire N2445;
wire N2446;
wire N2447;
wire N2448;
wire N2449;
wire N2450;
wire N2451;
wire N2452;
wire N2453;
wire N2454;
wire N2455;
wire N2456;
wire N2457;
wire N2458;
wire N2459;
wire N2460;
wire N2461;
wire N2462;
wire N2463;
wire N2464;
wire N2465;
wire N25;
wire N2500;
wire N2504;
wire N256;
wire N2570;
wire N2571;
wire N2572;
wire N2573;
wire N2574;
wire N2575;
wire N2576;
wire N2577;
wire N2593;
wire N2598;
wire N26;
wire N2607;
wire N2610;
wire N2613;
wire N2616;
wire N2619;
wire N2622;
wire N2625;
wire N2628;
wire N265;
wire N269;
wire N2696;
wire N27;
wire N2705;
wire N2709;
wire N2711;
wire N2713;
wire N2715;
wire N2717;
wire N2719;
wire N2721;
wire N2723;
wire N2724;
wire N2725;
wire N2726;
wire N2729;
wire N2732;
wire N2734;
wire N2736;
wire N2740;
wire N2744;
wire N2748;
wire N2752;
wire N2756;
wire N2760;
wire N2764;
wire N28;
wire N2837;
wire N2838;
wire N2847;
wire N285;
wire N2856;
wire N2857;
wire N2859;
wire N286;
wire N2861;
wire N2862;
wire N2863;
wire N2864;
wire N2865;
wire N2866;
wire N2867;
wire N2868;
wire N2869;
wire N287;
wire N2870;
wire N2871;
wire N2872;
wire N2873;
wire N2874;
wire N2875;
wire N2876;
wire N2877;
wire N2878;
wire N2879;
wire N2880;
wire N2881;
wire N2882;
wire N2883;
wire N2884;
wire N2885;
wire N2887;
wire N2888;
wire N2889;
wire N2890;
wire N2891;
wire N2892;
wire N2894;
wire N2929;
wire N2933;
wire N2993;
wire N2999;
wire N3000;
wire N3001;
wire N3002;
wire N3003;
wire N3004;
wire N3005;
wire N3006;
wire N3011;
wire N3020;
wire N3023;
wire N3033;
wire N3036;
wire N3039;
wire N3042;
wire N3045;
wire N3048;
wire N3051;
wire N3054;
wire N31;
wire N3124;
wire N3133;
wire N3134;
wire N3136;
wire N3138;
wire N3140;
wire N3142;
wire N3144;
wire N3146;
wire N3148;
wire N3150;
wire N3151;
wire N3153;
wire N3154;
wire N3156;
wire N3157;
wire N3158;
wire N3160;
wire N3164;
wire N3166;
wire N3168;
wire N317;
wire N3170;
wire N3174;
wire N3178;
wire N318;
wire N3182;
wire N3186;
wire N319;
wire N3190;
wire N3194;
wire N3198;
wire N32;
wire N320;
wire N321;
wire N322;
wire N323;
wire N3237;
wire N3238;
wire N324;
wire N325;
wire N326;
wire N327;
wire N3270;
wire N3271;
wire N3272;
wire N328;
wire N3289;
wire N329;
wire N3291;
wire N3292;
wire N3293;
wire N3294;
wire N3295;
wire N3296;
wire N3297;
wire N3298;
wire N3299;
wire N33;
wire N330;
wire N3300;
wire N3301;
wire N3302;
wire N3303;
wire N3304;
wire N3305;
wire N3306;
wire N3307;
wire N3308;
wire N3309;
wire N331;
wire N3310;
wire N3311;
wire N3312;
wire N3313;
wire N3314;
wire N3315;
wire N3316;
wire N3317;
wire N3318;
wire N3319;
wire N332;
wire N3320;
wire N3321;
wire N3322;
wire N3323;
wire N333;
wire N334;
wire N335;
wire N3358;
wire N3362;
wire N338;
wire N34;
wire N3428;
wire N3429;
wire N343;
wire N3430;
wire N3431;
wire N3432;
wire N3433;
wire N3434;
wire N3435;
wire N3450;
wire N3455;
wire N3464;
wire N3467;
wire N347;
wire N3470;
wire N3473;
wire N3476;
wire N3479;
wire N3482;
wire N3485;
wire N35;
wire N350;
wire N3554;
wire N3563;
wire N3565;
wire N3567;
wire N3569;
wire N3571;
wire N3573;
wire N3575;
wire N3577;
wire N3579;
wire N3580;
wire N3582;
wire N3583;
wire N3584;
wire N3585;
wire N3587;
wire N3590;
wire N3592;
wire N3594;
wire N3596;
wire N36;
wire N3600;
wire N3604;
wire N3608;
wire N3612;
wire N3616;
wire N3620;
wire N3624;
wire N364;
wire N3664;
wire N3665;
wire N3697;
wire N3698;
wire N3699;
wire N37;
wire N3716;
wire N3718;
wire N3719;
wire N372;
wire N3720;
wire N3721;
wire N3722;
wire N3723;
wire N3724;
wire N3725;
wire N3726;
wire N3727;
wire N3728;
wire N3729;
wire N3730;
wire N3731;
wire N3732;
wire N3733;
wire N3734;
wire N3735;
wire N3736;
wire N3737;
wire N3738;
wire N3739;
wire N3740;
wire N3741;
wire N3742;
wire N3743;
wire N3744;
wire N3745;
wire N3746;
wire N3747;
wire N3748;
wire N3749;
wire N3750;
wire N3785;
wire N3789;
wire N38;
wire N384;
wire N3856;
wire N3857;
wire N3858;
wire N3859;
wire N3860;
wire N3861;
wire N3862;
wire N3863;
wire N3878;
wire N3883;
wire N3892;
wire N3895;
wire N3898;
wire N39;
wire N390;
wire N3901;
wire N3904;
wire N3907;
wire N3910;
wire N3913;
wire N397;
wire N398;
wire N3982;
wire N399;
wire N3992;
wire N3994;
wire N3996;
wire N3998;
wire N40;
wire N4000;
wire N4002;
wire N4004;
wire N4006;
wire N4007;
wire N4009;
wire N4010;
wire N4011;
wire N4012;
wire N4014;
wire N4017;
wire N4019;
wire N4021;
wire N4025;
wire N4029;
wire N4033;
wire N4037;
wire N4041;
wire N4045;
wire N4049;
wire N4090;
wire N4091;
wire N4123;
wire N4124;
wire N4125;
wire N4142;
wire N4144;
wire N4145;
wire N4146;
wire N4147;
wire N4148;
wire N4149;
wire N4150;
wire N4151;
wire N4152;
wire N4153;
wire N4154;
wire N4155;
wire N4156;
wire N4157;
wire N4158;
wire N4159;
wire N4160;
wire N4161;
wire N4162;
wire N4163;
wire N4164;
wire N4165;
wire N4166;
wire N4167;
wire N4168;
wire N4169;
wire N4170;
wire N4171;
wire N4172;
wire N4173;
wire N4174;
wire N4175;
wire N4176;
wire N4211;
wire N4215;
wire N4281;
wire N4282;
wire N4283;
wire N4284;
wire N4285;
wire N4286;
wire N4287;
wire N4288;
wire N430;
wire N4303;
wire N4307;
wire N431;
wire N4316;
wire N4319;
wire N432;
wire N4322;
wire N4325;
wire N4328;
wire N433;
wire N4331;
wire N4334;
wire N4337;
wire N434;
wire N435;
wire N436;
wire N437;
wire N438;
wire N439;
wire N440;
wire N441;
wire N442;
wire N443;
wire N444;
wire N445;
wire N446;
wire N447;
wire N448;
wire N449;
wire N450;
wire N451;
wire N452;
wire N453;
wire N454;
wire N455;
wire N456;
wire N457;
wire N459;
wire N462;
wire N464;
wire N466;
wire N468;
wire N470;
wire N472;
wire N473;
wire N475;
wire N476;
wire N478;
wire N479;
wire N481;
wire N483;
wire N486;
wire N488;
wire N490;
wire N492;
wire N493;
wire N496;
wire N498;
wire N50;
wire N507;
wire N510;
wire N514;
wire N518;
wire N522;
wire N526;
wire N530;
wire N533;
wire N541;
wire N542;
wire N543;
wire N544;
wire N545;
wire N546;
wire N547;
wire N578;
wire N579;
wire N580;
wire N581;
wire N582;
wire N583;
wire N584;
wire N585;
wire N586;
wire N587;
wire N588;
wire N589;
wire N590;
wire N591;
wire N592;
wire N594;
wire N595;
wire N596;
wire N597;
wire N598;
wire N599;
wire N600;
wire N601;
wire N602;
wire N603;
wire N604;
wire N628;
wire N632;
wire N638;
wire N641;
wire N644;
wire N647;
wire N650;
wire N653;
wire N656;
wire N659;
wire N662;
wire N664;
wire N666;
wire N701;
wire N702;
wire N703;
wire N704;
wire N705;
wire N706;
wire N707;
wire N708;
wire N709;
wire N710;
wire N711;
wire N712;
wire N713;
wire N714;
wire N715;
wire N716;
wire N717;
wire N718;
wire N719;
wire N720;
wire N721;
wire N722;
wire N723;
wire N724;
wire N725;
wire N737;
wire N772;
wire N792;
wire N799;
wire N800;
wire N801;
wire N802;
wire N803;
wire N804;
wire N805;
wire N806;
wire N807;
wire N808;
wire N809;
wire N818;
wire N819;
wire N823;
wire N824;
wire N825;
wire N827;
wire N828;
wire N829;
wire N830;
wire N831;
wire N832;
wire N833;
wire N834;
wire N835;
wire N839;
wire N84;
wire N899;
wire N900;
wire N901;
wire N902;
wire N903;
wire N905;
wire N907;
wire N909;
wire N911;
wire N913;
wire N915;
wire N917;
wire N919;
wire N920;
wire N921;
wire N922;
wire N923;
wire N924;
wire N926;
wire N932;
wire N936;
wire N940;
wire N944;
wire N948;
wire N952;
wire N956;
wire N960;
wire N967;
wire N974;
nor #5 GDRQ(DRQ,N321);
nor #5 GHD0OUT(HD0OUT,N4007,N4012,N4142,N4175,N4215);
nor #5 GHD1OUT(HD1OUT,N3580,N3585,N3716,N3749,N3789);
nor #5 GHD2OUT(HD2OUT,N3151,N3158,N3289,N3322,N3362);
nor #5 GHD3OUT(HD3OUT,N2725,N2726,N2856,N2857,N2933);
nor #5 GHD4OUT(HD4OUT,N2296,N2301,N2432,N2464,N2504);
nor #5 GHD5OUT(HD5OUT,N1873,N1877,N2007,N2039,N2079);
nor #5 GHD6OUT(HD6OUT,N1335,N1336,N1436,N1437,N1458,N1588,N1620,N1687);
nor #5 GHD7OUT(HD7OUT,N1035,N1083,N1125,N1155,N1187,N899,N921,N967);
nor #5 GHDOEA(HDOEA,HCS,N116,N50);
nor #5 GHIRQ(HIRQ,N1432);
nor #5 GN1003(N1003,N903);
nor #5 GN1035(N1035,N1004,N441);
nor #5 GN1036(N1036,N1057,N459);
nor #5 GN1056(N1056,N34,N709);
nor #5 GN1083(N1083,N37,N664);
nor #5 GN1087(N1087,N120,N628);
nor #5 GN1125(N1125,N498,N919);
nor #5 GN1126(N1126,N1058,N442);
nor #5 GN115(N115,N124,N35);
nor #5 GN1155(N1155,N343,N84);
nor #5 GN116(N116,HO2);
nor #5 GN117(N117,N122);
nor #5 GN118(N118,N24);
nor #5 GN1187(N1187,N1082,N334);
nor #5 GN1188(N1188,N118,N1208);
nor #5 GN119(N119,N36);
nor #5 GN120(N120,N123);
nor #5 GN1206(N1206,N332,N595);
nor #5 GN1208(N1208,N321);
nor #5 GN121(N121,HCS,N116,N50);
nor #5 GN122(N122,HA0,HA2,N39);
nor #5 GN123(N123,N23,N32,PA0,PA2);
nor #5 GN124(N124,PCS,PNWDS);
nor #5 GN125(N125,N126,N176);
nor #5 GN126(N126,PCS,PNRDS);
nor #5 GN127(N127,N121);
nor #5 GN1314(N1314,N664);
nor #5 GN1326(N1326,N1346);
nor #5 GN1327(N1327,N708);
nor #5 GN1328(N1328,N1314,N34);
nor #5 GN1329(N1329,N118,N1339);
nor #5 GN1332(N1332,N1343,N321);
nor #5 GN1335(N1335,N318,N84);
nor #5 GN1336(N1336,N1327,N335);
nor #5 GN1339(N1339,N343);
nor #5 GN1343(N1343,N1434);
nor #5 GN1346(N1346,N4011,N4017,N4123);
nor #5 GN1398(N1398,N120,N1430);
nor #5 GN1399(N1399,N628);
nor #5 GN140(N140,N23,PA0,PA1,PA2);
nor #5 GN141(N141,HA0,HA1,HA2);
nor #5 GN1430(N1430,N666);
nor #5 GN1432(N1432,N1314,N1326);
nor #5 GN1433(N1433,N1876,N1882,N1988);
nor #5 GN1434(N1434,N2724,N2732,N2837);
nor #5 GN1435(N1435,N1349,N442);
nor #5 GN1436(N1436,N117,N1399);
nor #5 GN1437(N1437,N1396,N498);
nor #5 GN1453(N1453,N709);
nor #5 GN1455(N1455,N325,N454);
nor #5 GN1457(N1457,N1466,N435);
nor #5 GN1458(N1458,N1453,N37);
nor #5 GN1464(N1464,N1571,N924);
nor #5 GN1466(N1466,N1206,N1570,N1571);
nor #5 GN1536(N1536,N1456,N326);
nor #5 GN1570(N1570,N1206,N924);
nor #5 GN1588(N1588,N1538,N441);
nor #5 GN1616(N1616,N1537,N327);
nor #5 GN1620(N1620,N1612,N496);
nor #5 GN1687(N1687,N1614,N334);
nor #5 GN1688(N1688,N1589,N459);
nor #5 GN175(N175,N124,N35);
nor #5 GN176(N176,DACK,PNWDS);
nor #5 GN177(N177,N175,N459);
nor #5 GN1873(N1873,N1433,N335);
nor #5 GN1874(N1874,N1433,N325);
nor #5 GN1876(N1876,N1433,N1884);
nor #5 GN1877(N1877,N1872,N498);
nor #5 GN1879(N1879,N1875,N326);
nor #5 GN1882(N1882,N1990,N924);
nor #5 GN1884(N1884,N1206,N1988,N1990);
nor #5 GN1988(N1988,N1206,N924);
nor #5 GN1989(N1989,N1955,N327);
nor #5 GN2007(N2007,N1956,N441);
nor #5 GN2008(N2008,N2010,N442);
nor #5 GN2039(N2039,N2033,N496);
nor #5 GN2040(N2040,N2009,N459);
nor #5 GN207(N207,N119,N498);
nor #5 GN2079(N2079,N2035,N334);
nor #5 GN208(N208,N119,N496);
nor #5 GN209(N209,N175,N327);
nor #5 GN210(N210,N235,N237);
nor #5 GN211(N211,N23,N31,PA1,PA2);
nor #5 GN212(N212,N23,N31,N32,PA2);
nor #5 GN213(N213,N31,N33,PA1);
nor #5 GN214(N214,N23,N31,N32,N33);
nor #5 GN215(N215,N175,N326);
nor #5 GN216(N216,N228,N230);
nor #5 GN217(N217,N216,N231);
nor #5 GN218(N218,N210,N234);
nor #5 GN219(N219,N119,N335);
nor #5 GN220(N220,HA2,N39,N40);
nor #5 GN221(N221,HA1,N38,N40);
nor #5 GN222(N222,N38,N39,N40);
nor #5 GN223(N223,HA1,HA2,N40);
nor #5 GN228(N228,N323,N329,N330);
nor #5 GN2296(N2296,N269,N335);
nor #5 GN2298(N2298,N269,N325);
nor #5 GN23(N23,DACK);
nor #5 GN230(N230,N269);
nor #5 GN2300(N2300,N2308,N269);
nor #5 GN2301(N2301,N2295,N498);
nor #5 GN2303(N2303,N2299,N326);
nor #5 GN2306(N2306,N2415,N924);
nor #5 GN2308(N2308,N1206,N2412,N2415);
nor #5 GN231(N231,N256,N269);
nor #5 GN234(N234,N269,N320);
nor #5 GN235(N235,N269);
nor #5 GN237(N237,N333,N347,N436);
nor #5 GN24(N24,N23,N33,PA0,PA1);
nor #5 GN2412(N2412,N1206,N924);
nor #5 GN2414(N2414,N2379,N327);
nor #5 GN2432(N2432,N2380,N441);
nor #5 GN2433(N2433,N2435,N442);
nor #5 GN2464(N2464,N2458,N496);
nor #5 GN2465(N2465,N2434,N459);
nor #5 GN25(N25,N23,N32,N33,PA0);
nor #5 GN2504(N2504,N2460,N334);
nor #5 GN256(N256,N330);
nor #5 GN26(N26,N36);
nor #5 GN269(N269,N2300,N2306,N2412);
nor #5 GN27(N27,HA0,N38,N39);
nor #5 GN2724(N2724,N1434,N2734);
nor #5 GN2725(N2725,N2723,N496);
nor #5 GN2726(N2726,N2705,N498);
nor #5 GN2732(N2732,N2838,N924);
nor #5 GN2734(N2734,N1206,N2837,N2838);
nor #5 GN28(N28,HA0,HA1,N38);
nor #5 GN2837(N2837,N1206,N924);
nor #5 GN285(N285,N175,N442);
nor #5 GN2856(N2856,N2847,N334);
nor #5 GN2857(N2857,N1434,N335);
nor #5 GN286(N286,N119,N334);
nor #5 GN287(N287,N119,N441);
nor #5 GN2887(N2887,N1434,N325);
nor #5 GN2894(N2894,N2859,N326);
nor #5 GN2933(N2933,N2883,N441);
nor #5 GN2993(N2993,N2890,N327);
nor #5 GN3011(N3011,N2861,N442);
nor #5 GN3023(N3023,N2889,N459);
nor #5 GN31(N31,PA0);
nor #5 GN3133(N3133,N3157,N3166,N3270);
nor #5 GN3134(N3134,N1327,N3590);
nor #5 GN3151(N3151,N3133,N335);
nor #5 GN3153(N3153,N3133,N325);
nor #5 GN3156(N3156,N1453,N3164);
nor #5 GN3157(N3157,N3133,N3168);
nor #5 GN3158(N3158,N3150,N498);
nor #5 GN3160(N3160,N3154,N326);
nor #5 GN3164(N3164,N3133);
nor #5 GN3166(N3166,N3272,N924);
nor #5 GN3168(N3168,N1206,N3270,N3272);
nor #5 GN317(N317,N372);
nor #5 GN319(N319,N218,N317,N343);
nor #5 GN32(N32,PA1);
nor #5 GN320(N320,N333);
nor #5 GN321(N321,N265,N319);
nor #5 GN322(N322,N125,N326);
nor #5 GN324(N324,N127,N317,N498);
nor #5 GN325(N325,N140);
nor #5 GN326(N326,N213,N23);
nor #5 GN327(N327,N214);
nor #5 GN3270(N3270,N1206,N924);
nor #5 GN3271(N3271,N3237,N327);
nor #5 GN328(N328,N338);
nor #5 GN3289(N3289,N3238,N441);
nor #5 GN329(N329,N328,N592,N594,N632);
nor #5 GN3291(N3291,N3293,N442);
nor #5 GN33(N33,PA2);
nor #5 GN330(N330,N329,N737);
nor #5 GN331(N331,N323);
nor #5 GN332(N332,HRST);
nor #5 GN3322(N3322,N3316,N496);
nor #5 GN3323(N3323,N3292,N459);
nor #5 GN333(N333,N317,N347,N772);
nor #5 GN334(N334,N220);
nor #5 GN335(N335,N141);
nor #5 GN3362(N3362,N3318,N334);
nor #5 GN338(N338,N323);
nor #5 GN34(N34,N25);
nor #5 GN343(N343,N319,N398);
nor #5 GN347(N347,N440,N597,N662,N712);
nor #5 GN35(N35,DACK,PNRDS);
nor #5 GN350(N350,N324,N384,N431);
nor #5 GN3563(N3563,N3584,N3592,N3697);
nor #5 GN3580(N3580,N335,N3563);
nor #5 GN3582(N3582,N325,N3563);
nor #5 GN3584(N3584,N3563,N3594);
nor #5 GN3585(N3585,N3579,N498);
nor #5 GN3587(N3587,N326,N3583);
nor #5 GN3590(N3590,N3563);
nor #5 GN3592(N3592,N3699,N924);
nor #5 GN3594(N3594,N1206,N3697,N3699);
nor #5 GN36(N36,HCS,HRW,N116);
nor #5 GN3697(N3697,N1206,N924);
nor #5 GN3698(N3698,N327,N3664);
nor #5 GN37(N37,N27);
nor #5 GN3716(N3716,N3665,N441);
nor #5 GN3718(N3718,N3720,N442);
nor #5 GN372(N372,N332,N435);
nor #5 GN3749(N3749,N3743,N496);
nor #5 GN3750(N3750,N3719,N459);
nor #5 GN3789(N3789,N334,N3745);
nor #5 GN38(N38,HA2);
nor #5 GN384(N384,N350,N437);
nor #5 GN39(N39,HA1);
nor #5 GN398(N398,N320,N399);
nor #5 GN399(N399,N436);
nor #5 GN40(N40,HA0);
nor #5 GN4007(N4007,N1346,N335);
nor #5 GN4009(N4009,N1346,N325);
nor #5 GN4011(N4011,N1346,N4019);
nor #5 GN4012(N4012,N4006,N498);
nor #5 GN4014(N4014,N326,N4010);
nor #5 GN4017(N4017,N4125,N924);
nor #5 GN4019(N4019,N1206,N4123,N4125);
nor #5 GN4123(N4123,N1206,N924);
nor #5 GN4124(N4124,N327,N4090);
nor #5 GN4142(N4142,N4091,N441);
nor #5 GN4144(N4144,N4146,N442);
nor #5 GN4175(N4175,N4169,N496);
nor #5 GN4176(N4176,N4145,N459);
nor #5 GN4215(N4215,N334,N4171);
nor #5 GN430(N430,N317);
nor #5 GN431(N431,N116,N430);
nor #5 GN434(N434,N256,N331);
nor #5 GN435(N435,N1457,N1464,N1570);
nor #5 GN436(N436,N490,N597);
nor #5 GN438(N438,N127,N441);
nor #5 GN440(N440,N390,N438);
nor #5 GN441(N441,N221);
nor #5 GN442(N442,N211);
nor #5 GN444(N444,N285,N433,N507);
nor #5 GN445(N445,N455,N468,N510,N591);
nor #5 GN446(N446,N470,N472,N514,N579);
nor #5 GN447(N447,N473,N475,N518,N581);
nor #5 GN448(N448,N476,N478,N522,N583);
nor #5 GN449(N449,N479,N481,N526,N585);
nor #5 GN450(N450,N456,N483,N530,N587);
nor #5 GN451(N451,N486,N488,N533,N589);
nor #5 GN453(N453,N219,N466);
nor #5 GN455(N455,N445,N507,N638,N701);
nor #5 GN456(N456,N450,N526,N653,N706);
nor #5 GN457(N457,N324,N350);
nor #5 GN459(N459,N212);
nor #5 GN466(N466,N453,N595,N596);
nor #5 GN472(N472,N446,N591,N641,N702);
nor #5 GN475(N475,N447,N514,N644,N703);
nor #5 GN478(N478,N448,N518,N647,N704);
nor #5 GN481(N481,N449,N522,N650,N705);
nor #5 GN488(N488,N451,N530,N656,N707);
nor #5 GN490(N490,N317,N347,N436);
nor #5 GN496(N496,N222);
nor #5 GN498(N498,N223);
nor #5 GN50(N50,HRW);
nor #5 GN507(N507,N444,N454,N455,N800);
nor #5 GN510(N510,N541);
nor #5 GN514(N514,N446,N475,N542,N802);
nor #5 GN518(N518,N447,N478,N543,N803);
nor #5 GN522(N522,N448,N481,N544,N804);
nor #5 GN526(N526,N449,N456,N545,N805);
nor #5 GN530(N530,N450,N488,N546,N806);
nor #5 GN533(N533,N451,N547,N602,N807);
nor #5 GN579(N579,N542);
nor #5 GN581(N581,N543);
nor #5 GN583(N583,N544);
nor #5 GN585(N585,N545);
nor #5 GN587(N587,N546);
nor #5 GN589(N589,N547);
nor #5 GN591(N591,N445,N472,N541,N801);
nor #5 GN592(N592,N322,N432);
nor #5 GN594(N594,N287,N329,N462);
nor #5 GN595(N595,N219,N710,N799);
nor #5 GN596(N596,N219,N716,N799);
nor #5 GN597(N597,N215,N347,N492);
nor #5 GN598(N598,N125,N442);
nor #5 GN599(N599,N125,N459);
nor #5 GN600(N600,N125,N327);
nor #5 GN601(N601,N454);
nor #5 GN602(N602,N457,N533,N659,N711);
nor #5 GN603(N603,N127,N334);
nor #5 GN604(N604,N127,N496);
nor #5 GN628(N628,N317,N599,N714);
nor #5 GN632(N632,N330);
nor #5 GN662(N662,N333);
nor #5 GN664(N664,N317,N604,N724);
nor #5 GN666(N666,N317,N603,N725);
nor #5 GN701(N701,N468);
nor #5 GN702(N702,N470);
nor #5 GN703(N703,N473);
nor #5 GN704(N704,N476);
nor #5 GN705(N705,N479);
nor #5 GN706(N706,N483);
nor #5 GN707(N707,N486);
nor #5 GN708(N708,N317,N598,N713);
nor #5 GN709(N709,N317,N600,N715);
nor #5 GN712(N712,N835);
nor #5 GN713(N713,N207,N708);
nor #5 GN714(N714,N286,N628);
nor #5 GN715(N715,N208,N709);
nor #5 GN716(N716,N710);
nor #5 GN724(N724,N209,N664);
nor #5 GN725(N725,N177,N666);
nor #5 GN737(N737,N317,N330,N592);
nor #5 GN772(N772,N333,N440);
nor #5 GN792(N792,N437);
nor #5 GN799(N799,N902);
nor #5 GN800(N800,N638);
nor #5 GN801(N801,N641);
nor #5 GN802(N802,N644);
nor #5 GN803(N803,N647);
nor #5 GN804(N804,N650);
nor #5 GN805(N805,N653);
nor #5 GN806(N806,N656);
nor #5 GN807(N807,N711);
nor #5 GN808(N808,N286);
nor #5 GN809(N809,N208);
nor #5 GN818(N818,N209);
nor #5 GN819(N819,N177);
nor #5 GN824(N824,N207);
nor #5 GN835(N835,N436);
nor #5 GN84(N84,N28);
nor #5 GN899(N899,N117,N666);
nor #5 GN900(N900,N326,N923);
nor #5 GN901(N901,N974);
nor #5 GN902(N902,N901);
nor #5 GN903(N903,N453);
nor #5 GN921(N921,N496,N920);
nor #5 GN922(N922,N325,N708);
nor #5 GN924(N924,N332,N596);
nor #5 GN926(N926,N1002,N327);
nor #5 GN967(N967,N335,N792);
nor #5 GN974(N974,N1003);
nor #5 GPD0OUT(PD0OUT,N4009,N4014,N4124,N4144,N4176);
nor #5 GPD1OUT(PD1OUT,N3582,N3587,N3698,N3718,N3750);
nor #5 GPD2OUT(PD2OUT,N3153,N3160,N3271,N3291,N3323);
nor #5 GPD3OUT(PD3OUT,N2887,N2894,N2993,N3011,N3023);
nor #5 GPD4OUT(PD4OUT,N2298,N2303,N2414,N2433,N2465);
nor #5 GPD5OUT(PD5OUT,N1874,N1879,N1989,N2008,N2040);
nor #5 GPD6OUT(PD6OUT,N1328,N1329,N1398,N1435,N1455,N1536,N1616,N1688);
nor #5 GPD7OUT(PD7OUT,N1036,N1056,N1087,N1126,N1188,N900,N922,N926);
nor #5 GPDOEA(PDOEA,DACK,PNWDS);
nor #5 GPDOEB(PDOEB,PCS,PNRDS);
nor #5 GPIRQ(PIRQ,N3134,N3156);
nor #5 GPNMI(PNMI,N1332);
nor #5 GPRST(PRST,N1433,N332);
d_latch d0(.NQ(N1057),.D(N710),.EN(N808));
d_latch d1(.NQ(N1002),.D(N710),.EN(N809));
d_latch d10(.Q(N1075),.D(N915),.EN(N587));
d_latch d100(.Q(N2291),.D(N2575),.EN(N706));
d_latch d101(.Q(N2293),.D(N2576),.EN(N707));
d_latch d102(.NQ(N2295),.D(N2577),.EN(N792));
d_latch d103(.Q(N2415),.D(HD4IN),.EN(N26));
d_latch d104(.NQ(N2434),.D(N2415),.EN(N808));
d_latch d105(.NQ(N2379),.D(N2415),.EN(N809));
d_latch d106(.NQ(N2299),.D(N2439),.EN(N632));
d_latch d107(.Q(N2439),.D(N2415),.EN(N338));
d_latch d108(.Q(N2440),.D(N2271),.EN(N601));
d_latch d109(.Q(N2442),.D(N2281),.EN(N510));
d_latch d11(.Q(N1077),.D(N917),.EN(N589));
d_latch d110(.Q(N2444),.D(N2283),.EN(N579));
d_latch d111(.Q(N2446),.D(N2285),.EN(N581));
d_latch d112(.Q(N2448),.D(N2287),.EN(N583));
d_latch d113(.Q(N2450),.D(N2289),.EN(N585));
d_latch d114(.Q(N2452),.D(N2291),.EN(N587));
d_latch d115(.Q(N2454),.D(N2293),.EN(N589));
d_latch d116(.Q(N2456),.D(N2271),.EN(N835));
d_latch d117(.NQ(N2380),.D(N2456),.EN(N662));
d_latch d118(.NQ(N2458),.D(N2271),.EN(N818));
d_latch d119(.NQ(N2435),.D(N2415),.EN(N824));
d_latch d12(.Q(N1079),.D(N823),.EN(N835));
d_latch d120(.NQ(N2460),.D(N2271),.EN(N819));
d_latch d121(.Q(N2570),.D(N2440),.EN(N800));
d_latch d122(.Q(N2571),.D(N2442),.EN(N801));
d_latch d123(.Q(N2572),.D(N2444),.EN(N802));
d_latch d124(.Q(N2573),.D(N2446),.EN(N803));
d_latch d125(.Q(N2574),.D(N2448),.EN(N804));
d_latch d126(.Q(N2575),.D(N2450),.EN(N805));
d_latch d127(.Q(N2576),.D(N2452),.EN(N806));
d_latch d128(.Q(N2577),.D(N2454),.EN(N807));
d_latch d129(.NQ(N2271),.D(PD4IN),.EN(N115));
d_latch d13(.NQ(N1004),.D(N1079),.EN(N662));
d_latch d130(.Q(N2709),.D(N2999),.EN(N701));
d_latch d131(.Q(N2711),.D(N3000),.EN(N702));
d_latch d132(.Q(N2713),.D(N3001),.EN(N703));
d_latch d133(.Q(N2715),.D(N3002),.EN(N704));
d_latch d134(.Q(N2717),.D(N3003),.EN(N705));
d_latch d135(.Q(N2719),.D(N3004),.EN(N706));
d_latch d136(.Q(N2721),.D(N3005),.EN(N707));
d_latch d137(.NQ(N2696),.D(PD3IN),.EN(N115));
d_latch d138(.NQ(N2705),.D(N3006),.EN(N792));
d_latch d139(.Q(N2838),.D(HD3IN),.EN(N26));
d_latch d14(.NQ(N920),.D(N823),.EN(N818));
d_latch d140(.NQ(N2889),.D(N2838),.EN(N808));
d_latch d141(.NQ(N2890),.D(N2838),.EN(N809));
d_latch d142(.NQ(N2859),.D(N2865),.EN(N632));
d_latch d143(.Q(N2865),.D(N2838),.EN(N338));
d_latch d144(.Q(N2866),.D(N2696),.EN(N601));
d_latch d145(.Q(N2868),.D(N2709),.EN(N510));
d_latch d146(.Q(N2870),.D(N2711),.EN(N579));
d_latch d147(.Q(N2872),.D(N2713),.EN(N581));
d_latch d148(.Q(N2874),.D(N2715),.EN(N583));
d_latch d149(.Q(N2876),.D(N2717),.EN(N585));
d_latch d15(.NQ(N1058),.D(N710),.EN(N824));
d_latch d150(.Q(N2878),.D(N2719),.EN(N587));
d_latch d151(.Q(N2880),.D(N2721),.EN(N589));
d_latch d152(.Q(N2882),.D(N2696),.EN(N835));
d_latch d153(.NQ(N2883),.D(N2882),.EN(N662));
d_latch d154(.NQ(N2723),.D(N2696),.EN(N818));
d_latch d155(.NQ(N2861),.D(N2838),.EN(N824));
d_latch d156(.NQ(N2847),.D(N2696),.EN(N819));
d_latch d157(.Q(N2999),.D(N2866),.EN(N800));
d_latch d158(.Q(N3000),.D(N2868),.EN(N801));
d_latch d159(.Q(N3001),.D(N2870),.EN(N802));
d_latch d16(.NQ(N1082),.D(N823),.EN(N819));
d_latch d160(.Q(N3002),.D(N2872),.EN(N803));
d_latch d161(.Q(N3003),.D(N2874),.EN(N804));
d_latch d162(.Q(N3004),.D(N2876),.EN(N805));
d_latch d163(.Q(N3005),.D(N2878),.EN(N806));
d_latch d164(.Q(N3006),.D(N2880),.EN(N807));
d_latch d165(.Q(N3136),.D(N3428),.EN(N701));
d_latch d166(.Q(N3138),.D(N3429),.EN(N702));
d_latch d167(.Q(N3140),.D(N3430),.EN(N703));
d_latch d168(.Q(N3142),.D(N3431),.EN(N704));
d_latch d169(.Q(N3144),.D(N3432),.EN(N705));
d_latch d17(.Q(N1194),.D(N1063),.EN(N800));
d_latch d170(.Q(N3146),.D(N3433),.EN(N706));
d_latch d171(.Q(N3148),.D(N3434),.EN(N707));
d_latch d172(.NQ(N3150),.D(N3435),.EN(N792));
d_latch d173(.Q(N3272),.D(HD2IN),.EN(N26));
d_latch d174(.NQ(N3292),.D(N3272),.EN(N808));
d_latch d175(.NQ(N3237),.D(N3272),.EN(N809));
d_latch d176(.NQ(N3154),.D(N3297),.EN(N632));
d_latch d177(.Q(N3297),.D(N3272),.EN(N338));
d_latch d178(.Q(N3298),.D(N3124),.EN(N601));
d_latch d179(.Q(N3300),.D(N3136),.EN(N510));
d_latch d18(.Q(N1195),.D(N1065),.EN(N801));
d_latch d180(.Q(N3302),.D(N3138),.EN(N579));
d_latch d181(.Q(N3304),.D(N3140),.EN(N581));
d_latch d182(.Q(N3306),.D(N3142),.EN(N583));
d_latch d183(.Q(N3308),.D(N3144),.EN(N585));
d_latch d184(.Q(N3310),.D(N3146),.EN(N587));
d_latch d185(.Q(N3312),.D(N3148),.EN(N589));
d_latch d186(.Q(N3314),.D(N3124),.EN(N835));
d_latch d187(.NQ(N3238),.D(N3314),.EN(N662));
d_latch d188(.NQ(N3316),.D(N3124),.EN(N818));
d_latch d189(.NQ(N3293),.D(N3272),.EN(N824));
d_latch d19(.Q(N1196),.D(N1067),.EN(N802));
d_latch d190(.NQ(N3318),.D(N3124),.EN(N819));
d_latch d191(.Q(N3428),.D(N3298),.EN(N800));
d_latch d192(.Q(N3429),.D(N3300),.EN(N801));
d_latch d193(.Q(N3430),.D(N3302),.EN(N802));
d_latch d194(.Q(N3431),.D(N3304),.EN(N803));
d_latch d195(.Q(N3432),.D(N3306),.EN(N804));
d_latch d196(.Q(N3433),.D(N3308),.EN(N805));
d_latch d197(.Q(N3434),.D(N3310),.EN(N806));
d_latch d198(.Q(N3435),.D(N3312),.EN(N807));
d_latch d199(.NQ(N3124),.D(PD2IN),.EN(N115));
d_latch d2(.NQ(N923),.D(N1062),.EN(N632));
d_latch d20(.Q(N1197),.D(N1069),.EN(N803));
d_latch d200(.Q(N3565),.D(N3856),.EN(N701));
d_latch d201(.Q(N3567),.D(N3857),.EN(N702));
d_latch d202(.Q(N3569),.D(N3858),.EN(N703));
d_latch d203(.Q(N3571),.D(N3859),.EN(N704));
d_latch d204(.Q(N3573),.D(N3860),.EN(N705));
d_latch d205(.Q(N3575),.D(N3861),.EN(N706));
d_latch d206(.Q(N3577),.D(N3862),.EN(N707));
d_latch d207(.NQ(N3579),.D(N3863),.EN(N792));
d_latch d208(.Q(N3699),.D(HD1IN),.EN(N26));
d_latch d209(.NQ(N3719),.D(N3699),.EN(N808));
d_latch d21(.Q(N1198),.D(N1071),.EN(N804));
d_latch d210(.NQ(N3664),.D(N3699),.EN(N809));
d_latch d211(.NQ(N3583),.D(N3724),.EN(N632));
d_latch d212(.Q(N3724),.D(N3699),.EN(N338));
d_latch d213(.Q(N3725),.D(N3554),.EN(N601));
d_latch d214(.Q(N3727),.D(N3565),.EN(N510));
d_latch d215(.Q(N3729),.D(N3567),.EN(N579));
d_latch d216(.Q(N3731),.D(N3569),.EN(N581));
d_latch d217(.Q(N3733),.D(N3571),.EN(N583));
d_latch d218(.Q(N3735),.D(N3573),.EN(N585));
d_latch d219(.Q(N3737),.D(N3575),.EN(N587));
d_latch d22(.Q(N1199),.D(N1073),.EN(N805));
d_latch d220(.Q(N3739),.D(N3577),.EN(N589));
d_latch d221(.Q(N3741),.D(N3554),.EN(N835));
d_latch d222(.NQ(N3665),.D(N3741),.EN(N662));
d_latch d223(.NQ(N3743),.D(N3554),.EN(N818));
d_latch d224(.NQ(N3720),.D(N3699),.EN(N824));
d_latch d225(.NQ(N3745),.D(N3554),.EN(N819));
d_latch d226(.Q(N3856),.D(N3725),.EN(N800));
d_latch d227(.Q(N3857),.D(N3727),.EN(N801));
d_latch d228(.Q(N3858),.D(N3729),.EN(N802));
d_latch d229(.Q(N3859),.D(N3731),.EN(N803));
d_latch d23(.Q(N1200),.D(N1075),.EN(N806));
d_latch d230(.Q(N3860),.D(N3733),.EN(N804));
d_latch d231(.Q(N3861),.D(N3735),.EN(N805));
d_latch d232(.Q(N3862),.D(N3737),.EN(N806));
d_latch d233(.Q(N3863),.D(N3739),.EN(N807));
d_latch d234(.NQ(N3554),.D(PD1IN),.EN(N115));
d_latch d235(.Q(N3992),.D(N4281),.EN(N701));
d_latch d236(.Q(N3994),.D(N4282),.EN(N702));
d_latch d237(.Q(N3996),.D(N4283),.EN(N703));
d_latch d238(.Q(N3998),.D(N4284),.EN(N704));
d_latch d239(.Q(N4000),.D(N4285),.EN(N705));
d_latch d24(.Q(N1201),.D(N1077),.EN(N807));
d_latch d240(.Q(N4002),.D(N4286),.EN(N706));
d_latch d241(.Q(N4004),.D(N4287),.EN(N707));
d_latch d242(.NQ(N4006),.D(N4288),.EN(N792));
d_latch d243(.Q(N4125),.D(HD0IN),.EN(N26));
d_latch d244(.NQ(N4145),.D(N4125),.EN(N808));
d_latch d245(.NQ(N4090),.D(N4125),.EN(N809));
d_latch d246(.NQ(N4010),.D(N4150),.EN(N632));
d_latch d247(.Q(N4150),.D(N4125),.EN(N338));
d_latch d248(.Q(N4151),.D(N3982),.EN(N601));
d_latch d249(.Q(N4153),.D(N3992),.EN(N510));
d_latch d25(.Q(N1439),.D(N1724),.EN(N701));
d_latch d250(.Q(N4155),.D(N3994),.EN(N579));
d_latch d251(.Q(N4157),.D(N3996),.EN(N581));
d_latch d252(.Q(N4159),.D(N3998),.EN(N583));
d_latch d253(.Q(N4161),.D(N4000),.EN(N585));
d_latch d254(.Q(N4163),.D(N4002),.EN(N587));
d_latch d255(.Q(N4165),.D(N4004),.EN(N589));
d_latch d256(.Q(N4167),.D(N3982),.EN(N835));
d_latch d257(.NQ(N4091),.D(N4167),.EN(N662));
d_latch d258(.NQ(N4169),.D(N3982),.EN(N818));
d_latch d259(.NQ(N4146),.D(N4125),.EN(N824));
d_latch d26(.Q(N1441),.D(N1725),.EN(N702));
d_latch d260(.NQ(N4171),.D(N3982),.EN(N819));
d_latch d261(.Q(N4281),.D(N4151),.EN(N800));
d_latch d262(.Q(N4282),.D(N4153),.EN(N801));
d_latch d263(.Q(N4283),.D(N4155),.EN(N802));
d_latch d264(.Q(N4284),.D(N4157),.EN(N803));
d_latch d265(.Q(N4285),.D(N4159),.EN(N804));
d_latch d266(.Q(N4286),.D(N4161),.EN(N805));
d_latch d267(.Q(N4287),.D(N4163),.EN(N806));
d_latch d268(.Q(N4288),.D(N4165),.EN(N807));
d_latch d269(.NQ(N3982),.D(PD0IN),.EN(N115));
d_latch d27(.Q(N1443),.D(N1726),.EN(N703));
d_latch d270(.Q(N710),.D(HD7IN),.EN(N26));
d_latch d271(.NQ(N823),.D(PD7IN),.EN(N115));
d_latch d272(.Q(N905),.D(N1194),.EN(N701));
d_latch d273(.Q(N907),.D(N1195),.EN(N702));
d_latch d274(.Q(N909),.D(N1196),.EN(N703));
d_latch d275(.Q(N911),.D(N1197),.EN(N704));
d_latch d276(.Q(N913),.D(N1198),.EN(N705));
d_latch d277(.Q(N915),.D(N1199),.EN(N706));
d_latch d278(.Q(N917),.D(N1200),.EN(N707));
d_latch d279(.NQ(N919),.D(N1201),.EN(N792));
d_latch d28(.Q(N1445),.D(N1727),.EN(N704));
d_latch d29(.Q(N1447),.D(N1728),.EN(N705));
d_latch d3(.Q(N1062),.D(N710),.EN(N338));
d_latch d30(.Q(N1449),.D(N1729),.EN(N706));
d_latch d31(.Q(N1451),.D(N1730),.EN(N707));
d_latch d32(.NQ(N1396),.D(N1731),.EN(N792));
d_latch d33(.Q(N1571),.D(HD6IN),.EN(N26));
d_latch d34(.NQ(N1589),.D(N1571),.EN(N808));
d_latch d35(.NQ(N1537),.D(N1571),.EN(N809));
d_latch d36(.NQ(N1456),.D(N1593),.EN(N632));
d_latch d37(.Q(N1593),.D(N1571),.EN(N338));
d_latch d38(.Q(N1594),.D(N1431),.EN(N601));
d_latch d39(.Q(N1596),.D(N1439),.EN(N510));
d_latch d4(.Q(N1063),.D(N823),.EN(N601));
d_latch d40(.Q(N1598),.D(N1441),.EN(N579));
d_latch d41(.Q(N1600),.D(N1443),.EN(N581));
d_latch d42(.Q(N1602),.D(N1445),.EN(N583));
d_latch d43(.Q(N1604),.D(N1447),.EN(N585));
d_latch d44(.Q(N1606),.D(N1449),.EN(N587));
d_latch d45(.Q(N1608),.D(N1451),.EN(N589));
d_latch d46(.Q(N1610),.D(N1431),.EN(N835));
d_latch d47(.NQ(N1538),.D(N1610),.EN(N662));
d_latch d48(.NQ(N1612),.D(N1431),.EN(N818));
d_latch d49(.NQ(N1349),.D(N1571),.EN(N824));
d_latch d5(.Q(N1065),.D(N905),.EN(N510));
d_latch d50(.NQ(N1614),.D(N1431),.EN(N819));
d_latch d51(.Q(N1724),.D(N1594),.EN(N800));
d_latch d52(.Q(N1725),.D(N1596),.EN(N801));
d_latch d53(.Q(N1726),.D(N1598),.EN(N802));
d_latch d54(.Q(N1727),.D(N1600),.EN(N803));
d_latch d55(.Q(N1728),.D(N1602),.EN(N804));
d_latch d56(.Q(N1729),.D(N1604),.EN(N805));
d_latch d57(.Q(N1730),.D(N1606),.EN(N806));
d_latch d58(.Q(N1731),.D(N1608),.EN(N807));
d_latch d59(.NQ(N1431),.D(PD6IN),.EN(N115));
d_latch d6(.Q(N1067),.D(N907),.EN(N579));
d_latch d60(.Q(N1858),.D(N2145),.EN(N701));
d_latch d61(.Q(N1860),.D(N2146),.EN(N702));
d_latch d62(.Q(N1862),.D(N2147),.EN(N703));
d_latch d63(.Q(N1864),.D(N2148),.EN(N704));
d_latch d64(.Q(N1866),.D(N2149),.EN(N705));
d_latch d65(.Q(N1868),.D(N2150),.EN(N706));
d_latch d66(.Q(N1870),.D(N2151),.EN(N707));
d_latch d67(.NQ(N1872),.D(N2152),.EN(N792));
d_latch d68(.Q(N1990),.D(HD5IN),.EN(N26));
d_latch d69(.NQ(N2009),.D(N1990),.EN(N808));
d_latch d7(.Q(N1069),.D(N909),.EN(N581));
d_latch d70(.NQ(N1955),.D(N1990),.EN(N809));
d_latch d71(.NQ(N1875),.D(N2014),.EN(N632));
d_latch d72(.Q(N2014),.D(N1990),.EN(N338));
d_latch d73(.Q(N2015),.D(N1848),.EN(N601));
d_latch d74(.Q(N2017),.D(N1858),.EN(N510));
d_latch d75(.Q(N2019),.D(N1860),.EN(N579));
d_latch d76(.Q(N2021),.D(N1862),.EN(N581));
d_latch d77(.Q(N2023),.D(N1864),.EN(N583));
d_latch d78(.Q(N2025),.D(N1866),.EN(N585));
d_latch d79(.Q(N2027),.D(N1868),.EN(N587));
d_latch d8(.Q(N1071),.D(N911),.EN(N583));
d_latch d80(.Q(N2029),.D(N1870),.EN(N589));
d_latch d81(.Q(N2031),.D(N1848),.EN(N835));
d_latch d82(.NQ(N1956),.D(N2031),.EN(N662));
d_latch d83(.NQ(N2033),.D(N1848),.EN(N818));
d_latch d84(.NQ(N2010),.D(N1990),.EN(N824));
d_latch d85(.NQ(N2035),.D(N1848),.EN(N819));
d_latch d86(.Q(N2145),.D(N2015),.EN(N800));
d_latch d87(.Q(N2146),.D(N2017),.EN(N801));
d_latch d88(.Q(N2147),.D(N2019),.EN(N802));
d_latch d89(.Q(N2148),.D(N2021),.EN(N803));
d_latch d9(.Q(N1073),.D(N913),.EN(N585));
d_latch d90(.Q(N2149),.D(N2023),.EN(N804));
d_latch d91(.Q(N2150),.D(N2025),.EN(N805));
d_latch d92(.Q(N2151),.D(N2027),.EN(N806));
d_latch d93(.Q(N2152),.D(N2029),.EN(N807));
d_latch d94(.NQ(N1848),.D(PD5IN),.EN(N115));
d_latch d95(.Q(N2281),.D(N2570),.EN(N701));
d_latch d96(.Q(N2283),.D(N2571),.EN(N702));
d_latch d97(.Q(N2285),.D(N2572),.EN(N703));
d_latch d98(.Q(N2287),.D(N2573),.EN(N704));
d_latch d99(.Q(N2289),.D(N2574),.EN(N705));
sr_latch sr0(.NQ(N318),.Q(N265),.R(N434),.S(N217));
sr_latch sr1(.NQ(N464),.Q(N323),.R(N594),.S(N329));
sr_latch sr10(.Q(N470),.R(N472),.S(N446));
sr_latch sr11(.Q(N473),.R(N475),.S(N447));
sr_latch sr12(.Q(N476),.R(N478),.S(N448));
sr_latch sr13(.Q(N479),.R(N481),.S(N449));
sr_latch sr14(.Q(N483),.R(N456),.S(N450));
sr_latch sr15(.Q(N486),.R(N488),.S(N451));
sr_latch sr16(.Q(N541),.R(N445),.S(N591));
sr_latch sr17(.Q(N542),.R(N446),.S(N514));
sr_latch sr18(.Q(N543),.R(N447),.S(N518));
sr_latch sr19(.Q(N544),.R(N448),.S(N522));
sr_latch sr2(.NQ(N454),.Q(N364),.R(N507),.S(N444));
sr_latch sr20(.Q(N545),.R(N449),.S(N526));
sr_latch sr21(.Q(N546),.R(N450),.S(N530));
sr_latch sr22(.Q(N547),.R(N451),.S(N533));
sr_latch sr23(.Q(N638),.R(N507),.S(N455));
sr_latch sr24(.Q(N641),.R(N591),.S(N472));
sr_latch sr25(.Q(N644),.R(N514),.S(N475));
sr_latch sr26(.Q(N647),.R(N518),.S(N478));
sr_latch sr27(.Q(N650),.R(N522),.S(N481));
sr_latch sr28(.Q(N653),.R(N526),.S(N456));
sr_latch sr29(.Q(N656),.R(N530),.S(N488));
sr_latch sr3(.Q(N390),.R(N438),.S(N333));
sr_latch sr30(.Q(N711),.R(N533),.S(N602));
sr_latch sr4(.NQ(N433),.R(N364),.S(N285));
sr_latch sr5(.Q(N432),.R(N322),.S(N330));
sr_latch sr6(.NQ(N659),.Q(N437),.R(N602),.S(N457));
sr_latch sr7(.NQ(N462),.R(N464),.S(N287));
sr_latch sr8(.NQ(N492),.R(N490),.S(N215));
sr_latch sr9(.Q(N468),.R(N455),.S(N445));
endmodule
